`include "/home/wzc/master_project/verilog/systolic_array/32bit_PE.v"
module SA64(rst, clk, weight_en, in_weight_0, in_psum_0, in_weight_1, in_psum_1, in_weight_2, in_psum_2, in_weight_3, in_psum_3, in_weight_4, in_psum_4, in_weight_5, in_psum_5, in_weight_6, in_psum_6, in_weight_7, in_psum_7, in_weight_8, in_psum_8, in_weight_9, in_psum_9, in_weight_10, in_psum_10, in_weight_11, in_psum_11, in_weight_12, in_psum_12, in_weight_13, in_psum_13, in_weight_14, in_psum_14, in_weight_15, in_psum_15, in_weight_16, in_psum_16, in_weight_17, in_psum_17, in_weight_18, in_psum_18, in_weight_19, in_psum_19, in_weight_20, in_psum_20, in_weight_21, in_psum_21, in_weight_22, in_psum_22, in_weight_23, in_psum_23, in_weight_24, in_psum_24, in_weight_25, in_psum_25, in_weight_26, in_psum_26, in_weight_27, in_psum_27, in_weight_28, in_psum_28, in_weight_29, in_psum_29, in_weight_30, in_psum_30, in_weight_31, in_psum_31, in_weight_32, in_psum_32, in_weight_33, in_psum_33, in_weight_34, in_psum_34, in_weight_35, in_psum_35, in_weight_36, in_psum_36, in_weight_37, in_psum_37, in_weight_38, in_psum_38, in_weight_39, in_psum_39, in_weight_40, in_psum_40, in_weight_41, in_psum_41, in_weight_42, in_psum_42, in_weight_43, in_psum_43, in_weight_44, in_psum_44, in_weight_45, in_psum_45, in_weight_46, in_psum_46, in_weight_47, in_psum_47, in_weight_48, in_psum_48, in_weight_49, in_psum_49, in_weight_50, in_psum_50, in_weight_51, in_psum_51, in_weight_52, in_psum_52, in_weight_53, in_psum_53, in_weight_54, in_psum_54, in_weight_55, in_psum_55, in_weight_56, in_psum_56, in_weight_57, in_psum_57, in_weight_58, in_psum_58, in_weight_59, in_psum_59, in_weight_60, in_psum_60, in_weight_61, in_psum_61, in_weight_62, in_psum_62, in_weight_63, in_psum_63, in_activation_0, in_activation_1, in_activation_2, in_activation_3, in_activation_4, in_activation_5, in_activation_6, in_activation_7, in_activation_8, in_activation_9, in_activation_10, in_activation_11, in_activation_12, in_activation_13, in_activation_14, in_activation_15, in_activation_16, in_activation_17, in_activation_18, in_activation_19, in_activation_20, in_activation_21, in_activation_22, in_activation_23, in_activation_24, in_activation_25, in_activation_26, in_activation_27, in_activation_28, in_activation_29, in_activation_30, in_activation_31, in_activation_32, in_activation_33, in_activation_34, in_activation_35, in_activation_36, in_activation_37, in_activation_38, in_activation_39, in_activation_40, in_activation_41, in_activation_42, in_activation_43, in_activation_44, in_activation_45, in_activation_46, in_activation_47, in_activation_48, in_activation_49, in_activation_50, in_activation_51, in_activation_52, in_activation_53, in_activation_54, in_activation_55, in_activation_56, in_activation_57, in_activation_58, in_activation_59, in_activation_60, in_activation_61, in_activation_62, in_activation_63, out_psum_0, out_psum_1, out_psum_2, out_psum_3, out_psum_4, out_psum_5, out_psum_6, out_psum_7, out_psum_8, out_psum_9, out_psum_10, out_psum_11, out_psum_12, out_psum_13, out_psum_14, out_psum_15, out_psum_16, out_psum_17, out_psum_18, out_psum_19, out_psum_20, out_psum_21, out_psum_22, out_psum_23, out_psum_24, out_psum_25, out_psum_26, out_psum_27, out_psum_28, out_psum_29, out_psum_30, out_psum_31, out_psum_32, out_psum_33, out_psum_34, out_psum_35, out_psum_36, out_psum_37, out_psum_38, out_psum_39, out_psum_40, out_psum_41, out_psum_42, out_psum_43, out_psum_44, out_psum_45, out_psum_46, out_psum_47, out_psum_48, out_psum_49, out_psum_50, out_psum_51, out_psum_52, out_psum_53, out_psum_54, out_psum_55, out_psum_56, out_psum_57, out_psum_58, out_psum_59, out_psum_60, out_psum_61, out_psum_62, out_psum_63);
input weight_en;
input clk,rst;
input signed[31:0]   in_weight_0;
input signed[31:0]   in_psum_0;
input signed[31:0]   in_weight_1;
input signed[31:0]   in_psum_1;
input signed[31:0]   in_weight_2;
input signed[31:0]   in_psum_2;
input signed[31:0]   in_weight_3;
input signed[31:0]   in_psum_3;
input signed[31:0]   in_weight_4;
input signed[31:0]   in_psum_4;
input signed[31:0]   in_weight_5;
input signed[31:0]   in_psum_5;
input signed[31:0]   in_weight_6;
input signed[31:0]   in_psum_6;
input signed[31:0]   in_weight_7;
input signed[31:0]   in_psum_7;
input signed[31:0]   in_weight_8;
input signed[31:0]   in_psum_8;
input signed[31:0]   in_weight_9;
input signed[31:0]   in_psum_9;
input signed[31:0]   in_weight_10;
input signed[31:0]   in_psum_10;
input signed[31:0]   in_weight_11;
input signed[31:0]   in_psum_11;
input signed[31:0]   in_weight_12;
input signed[31:0]   in_psum_12;
input signed[31:0]   in_weight_13;
input signed[31:0]   in_psum_13;
input signed[31:0]   in_weight_14;
input signed[31:0]   in_psum_14;
input signed[31:0]   in_weight_15;
input signed[31:0]   in_psum_15;
input signed[31:0]   in_weight_16;
input signed[31:0]   in_psum_16;
input signed[31:0]   in_weight_17;
input signed[31:0]   in_psum_17;
input signed[31:0]   in_weight_18;
input signed[31:0]   in_psum_18;
input signed[31:0]   in_weight_19;
input signed[31:0]   in_psum_19;
input signed[31:0]   in_weight_20;
input signed[31:0]   in_psum_20;
input signed[31:0]   in_weight_21;
input signed[31:0]   in_psum_21;
input signed[31:0]   in_weight_22;
input signed[31:0]   in_psum_22;
input signed[31:0]   in_weight_23;
input signed[31:0]   in_psum_23;
input signed[31:0]   in_weight_24;
input signed[31:0]   in_psum_24;
input signed[31:0]   in_weight_25;
input signed[31:0]   in_psum_25;
input signed[31:0]   in_weight_26;
input signed[31:0]   in_psum_26;
input signed[31:0]   in_weight_27;
input signed[31:0]   in_psum_27;
input signed[31:0]   in_weight_28;
input signed[31:0]   in_psum_28;
input signed[31:0]   in_weight_29;
input signed[31:0]   in_psum_29;
input signed[31:0]   in_weight_30;
input signed[31:0]   in_psum_30;
input signed[31:0]   in_weight_31;
input signed[31:0]   in_psum_31;
input signed[31:0]   in_weight_32;
input signed[31:0]   in_psum_32;
input signed[31:0]   in_weight_33;
input signed[31:0]   in_psum_33;
input signed[31:0]   in_weight_34;
input signed[31:0]   in_psum_34;
input signed[31:0]   in_weight_35;
input signed[31:0]   in_psum_35;
input signed[31:0]   in_weight_36;
input signed[31:0]   in_psum_36;
input signed[31:0]   in_weight_37;
input signed[31:0]   in_psum_37;
input signed[31:0]   in_weight_38;
input signed[31:0]   in_psum_38;
input signed[31:0]   in_weight_39;
input signed[31:0]   in_psum_39;
input signed[31:0]   in_weight_40;
input signed[31:0]   in_psum_40;
input signed[31:0]   in_weight_41;
input signed[31:0]   in_psum_41;
input signed[31:0]   in_weight_42;
input signed[31:0]   in_psum_42;
input signed[31:0]   in_weight_43;
input signed[31:0]   in_psum_43;
input signed[31:0]   in_weight_44;
input signed[31:0]   in_psum_44;
input signed[31:0]   in_weight_45;
input signed[31:0]   in_psum_45;
input signed[31:0]   in_weight_46;
input signed[31:0]   in_psum_46;
input signed[31:0]   in_weight_47;
input signed[31:0]   in_psum_47;
input signed[31:0]   in_weight_48;
input signed[31:0]   in_psum_48;
input signed[31:0]   in_weight_49;
input signed[31:0]   in_psum_49;
input signed[31:0]   in_weight_50;
input signed[31:0]   in_psum_50;
input signed[31:0]   in_weight_51;
input signed[31:0]   in_psum_51;
input signed[31:0]   in_weight_52;
input signed[31:0]   in_psum_52;
input signed[31:0]   in_weight_53;
input signed[31:0]   in_psum_53;
input signed[31:0]   in_weight_54;
input signed[31:0]   in_psum_54;
input signed[31:0]   in_weight_55;
input signed[31:0]   in_psum_55;
input signed[31:0]   in_weight_56;
input signed[31:0]   in_psum_56;
input signed[31:0]   in_weight_57;
input signed[31:0]   in_psum_57;
input signed[31:0]   in_weight_58;
input signed[31:0]   in_psum_58;
input signed[31:0]   in_weight_59;
input signed[31:0]   in_psum_59;
input signed[31:0]   in_weight_60;
input signed[31:0]   in_psum_60;
input signed[31:0]   in_weight_61;
input signed[31:0]   in_psum_61;
input signed[31:0]   in_weight_62;
input signed[31:0]   in_psum_62;
input signed[31:0]   in_weight_63;
input signed[31:0]   in_psum_63;
input signed[31:0]   in_activation_0;
input signed[31:0]   in_activation_1;
input signed[31:0]   in_activation_2;
input signed[31:0]   in_activation_3;
input signed[31:0]   in_activation_4;
input signed[31:0]   in_activation_5;
input signed[31:0]   in_activation_6;
input signed[31:0]   in_activation_7;
input signed[31:0]   in_activation_8;
input signed[31:0]   in_activation_9;
input signed[31:0]   in_activation_10;
input signed[31:0]   in_activation_11;
input signed[31:0]   in_activation_12;
input signed[31:0]   in_activation_13;
input signed[31:0]   in_activation_14;
input signed[31:0]   in_activation_15;
input signed[31:0]   in_activation_16;
input signed[31:0]   in_activation_17;
input signed[31:0]   in_activation_18;
input signed[31:0]   in_activation_19;
input signed[31:0]   in_activation_20;
input signed[31:0]   in_activation_21;
input signed[31:0]   in_activation_22;
input signed[31:0]   in_activation_23;
input signed[31:0]   in_activation_24;
input signed[31:0]   in_activation_25;
input signed[31:0]   in_activation_26;
input signed[31:0]   in_activation_27;
input signed[31:0]   in_activation_28;
input signed[31:0]   in_activation_29;
input signed[31:0]   in_activation_30;
input signed[31:0]   in_activation_31;
input signed[31:0]   in_activation_32;
input signed[31:0]   in_activation_33;
input signed[31:0]   in_activation_34;
input signed[31:0]   in_activation_35;
input signed[31:0]   in_activation_36;
input signed[31:0]   in_activation_37;
input signed[31:0]   in_activation_38;
input signed[31:0]   in_activation_39;
input signed[31:0]   in_activation_40;
input signed[31:0]   in_activation_41;
input signed[31:0]   in_activation_42;
input signed[31:0]   in_activation_43;
input signed[31:0]   in_activation_44;
input signed[31:0]   in_activation_45;
input signed[31:0]   in_activation_46;
input signed[31:0]   in_activation_47;
input signed[31:0]   in_activation_48;
input signed[31:0]   in_activation_49;
input signed[31:0]   in_activation_50;
input signed[31:0]   in_activation_51;
input signed[31:0]   in_activation_52;
input signed[31:0]   in_activation_53;
input signed[31:0]   in_activation_54;
input signed[31:0]   in_activation_55;
input signed[31:0]   in_activation_56;
input signed[31:0]   in_activation_57;
input signed[31:0]   in_activation_58;
input signed[31:0]   in_activation_59;
input signed[31:0]   in_activation_60;
input signed[31:0]   in_activation_61;
input signed[31:0]   in_activation_62;
input signed[31:0]   in_activation_63;
output signed[31:0]   out_psum_0;
output signed[31:0]   out_psum_1;
output signed[31:0]   out_psum_2;
output signed[31:0]   out_psum_3;
output signed[31:0]   out_psum_4;
output signed[31:0]   out_psum_5;
output signed[31:0]   out_psum_6;
output signed[31:0]   out_psum_7;
output signed[31:0]   out_psum_8;
output signed[31:0]   out_psum_9;
output signed[31:0]   out_psum_10;
output signed[31:0]   out_psum_11;
output signed[31:0]   out_psum_12;
output signed[31:0]   out_psum_13;
output signed[31:0]   out_psum_14;
output signed[31:0]   out_psum_15;
output signed[31:0]   out_psum_16;
output signed[31:0]   out_psum_17;
output signed[31:0]   out_psum_18;
output signed[31:0]   out_psum_19;
output signed[31:0]   out_psum_20;
output signed[31:0]   out_psum_21;
output signed[31:0]   out_psum_22;
output signed[31:0]   out_psum_23;
output signed[31:0]   out_psum_24;
output signed[31:0]   out_psum_25;
output signed[31:0]   out_psum_26;
output signed[31:0]   out_psum_27;
output signed[31:0]   out_psum_28;
output signed[31:0]   out_psum_29;
output signed[31:0]   out_psum_30;
output signed[31:0]   out_psum_31;
output signed[31:0]   out_psum_32;
output signed[31:0]   out_psum_33;
output signed[31:0]   out_psum_34;
output signed[31:0]   out_psum_35;
output signed[31:0]   out_psum_36;
output signed[31:0]   out_psum_37;
output signed[31:0]   out_psum_38;
output signed[31:0]   out_psum_39;
output signed[31:0]   out_psum_40;
output signed[31:0]   out_psum_41;
output signed[31:0]   out_psum_42;
output signed[31:0]   out_psum_43;
output signed[31:0]   out_psum_44;
output signed[31:0]   out_psum_45;
output signed[31:0]   out_psum_46;
output signed[31:0]   out_psum_47;
output signed[31:0]   out_psum_48;
output signed[31:0]   out_psum_49;
output signed[31:0]   out_psum_50;
output signed[31:0]   out_psum_51;
output signed[31:0]   out_psum_52;
output signed[31:0]   out_psum_53;
output signed[31:0]   out_psum_54;
output signed[31:0]   out_psum_55;
output signed[31:0]   out_psum_56;
output signed[31:0]   out_psum_57;
output signed[31:0]   out_psum_58;
output signed[31:0]   out_psum_59;
output signed[31:0]   out_psum_60;
output signed[31:0]   out_psum_61;
output signed[31:0]   out_psum_62;
output signed[31:0]   out_psum_63;
wire signed[31:0]    reg_activation_0_0;
wire signed[31:0]    reg_activation_0_1;
wire signed[31:0]    reg_activation_0_2;
wire signed[31:0]    reg_activation_0_3;
wire signed[31:0]    reg_activation_0_4;
wire signed[31:0]    reg_activation_0_5;
wire signed[31:0]    reg_activation_0_6;
wire signed[31:0]    reg_activation_0_7;
wire signed[31:0]    reg_activation_0_8;
wire signed[31:0]    reg_activation_0_9;
wire signed[31:0]    reg_activation_0_10;
wire signed[31:0]    reg_activation_0_11;
wire signed[31:0]    reg_activation_0_12;
wire signed[31:0]    reg_activation_0_13;
wire signed[31:0]    reg_activation_0_14;
wire signed[31:0]    reg_activation_0_15;
wire signed[31:0]    reg_activation_0_16;
wire signed[31:0]    reg_activation_0_17;
wire signed[31:0]    reg_activation_0_18;
wire signed[31:0]    reg_activation_0_19;
wire signed[31:0]    reg_activation_0_20;
wire signed[31:0]    reg_activation_0_21;
wire signed[31:0]    reg_activation_0_22;
wire signed[31:0]    reg_activation_0_23;
wire signed[31:0]    reg_activation_0_24;
wire signed[31:0]    reg_activation_0_25;
wire signed[31:0]    reg_activation_0_26;
wire signed[31:0]    reg_activation_0_27;
wire signed[31:0]    reg_activation_0_28;
wire signed[31:0]    reg_activation_0_29;
wire signed[31:0]    reg_activation_0_30;
wire signed[31:0]    reg_activation_0_31;
wire signed[31:0]    reg_activation_0_32;
wire signed[31:0]    reg_activation_0_33;
wire signed[31:0]    reg_activation_0_34;
wire signed[31:0]    reg_activation_0_35;
wire signed[31:0]    reg_activation_0_36;
wire signed[31:0]    reg_activation_0_37;
wire signed[31:0]    reg_activation_0_38;
wire signed[31:0]    reg_activation_0_39;
wire signed[31:0]    reg_activation_0_40;
wire signed[31:0]    reg_activation_0_41;
wire signed[31:0]    reg_activation_0_42;
wire signed[31:0]    reg_activation_0_43;
wire signed[31:0]    reg_activation_0_44;
wire signed[31:0]    reg_activation_0_45;
wire signed[31:0]    reg_activation_0_46;
wire signed[31:0]    reg_activation_0_47;
wire signed[31:0]    reg_activation_0_48;
wire signed[31:0]    reg_activation_0_49;
wire signed[31:0]    reg_activation_0_50;
wire signed[31:0]    reg_activation_0_51;
wire signed[31:0]    reg_activation_0_52;
wire signed[31:0]    reg_activation_0_53;
wire signed[31:0]    reg_activation_0_54;
wire signed[31:0]    reg_activation_0_55;
wire signed[31:0]    reg_activation_0_56;
wire signed[31:0]    reg_activation_0_57;
wire signed[31:0]    reg_activation_0_58;
wire signed[31:0]    reg_activation_0_59;
wire signed[31:0]    reg_activation_0_60;
wire signed[31:0]    reg_activation_0_61;
wire signed[31:0]    reg_activation_0_62;
wire signed[31:0]    reg_activation_0_63;
wire signed[31:0]    reg_activation_1_0;
wire signed[31:0]    reg_activation_1_1;
wire signed[31:0]    reg_activation_1_2;
wire signed[31:0]    reg_activation_1_3;
wire signed[31:0]    reg_activation_1_4;
wire signed[31:0]    reg_activation_1_5;
wire signed[31:0]    reg_activation_1_6;
wire signed[31:0]    reg_activation_1_7;
wire signed[31:0]    reg_activation_1_8;
wire signed[31:0]    reg_activation_1_9;
wire signed[31:0]    reg_activation_1_10;
wire signed[31:0]    reg_activation_1_11;
wire signed[31:0]    reg_activation_1_12;
wire signed[31:0]    reg_activation_1_13;
wire signed[31:0]    reg_activation_1_14;
wire signed[31:0]    reg_activation_1_15;
wire signed[31:0]    reg_activation_1_16;
wire signed[31:0]    reg_activation_1_17;
wire signed[31:0]    reg_activation_1_18;
wire signed[31:0]    reg_activation_1_19;
wire signed[31:0]    reg_activation_1_20;
wire signed[31:0]    reg_activation_1_21;
wire signed[31:0]    reg_activation_1_22;
wire signed[31:0]    reg_activation_1_23;
wire signed[31:0]    reg_activation_1_24;
wire signed[31:0]    reg_activation_1_25;
wire signed[31:0]    reg_activation_1_26;
wire signed[31:0]    reg_activation_1_27;
wire signed[31:0]    reg_activation_1_28;
wire signed[31:0]    reg_activation_1_29;
wire signed[31:0]    reg_activation_1_30;
wire signed[31:0]    reg_activation_1_31;
wire signed[31:0]    reg_activation_1_32;
wire signed[31:0]    reg_activation_1_33;
wire signed[31:0]    reg_activation_1_34;
wire signed[31:0]    reg_activation_1_35;
wire signed[31:0]    reg_activation_1_36;
wire signed[31:0]    reg_activation_1_37;
wire signed[31:0]    reg_activation_1_38;
wire signed[31:0]    reg_activation_1_39;
wire signed[31:0]    reg_activation_1_40;
wire signed[31:0]    reg_activation_1_41;
wire signed[31:0]    reg_activation_1_42;
wire signed[31:0]    reg_activation_1_43;
wire signed[31:0]    reg_activation_1_44;
wire signed[31:0]    reg_activation_1_45;
wire signed[31:0]    reg_activation_1_46;
wire signed[31:0]    reg_activation_1_47;
wire signed[31:0]    reg_activation_1_48;
wire signed[31:0]    reg_activation_1_49;
wire signed[31:0]    reg_activation_1_50;
wire signed[31:0]    reg_activation_1_51;
wire signed[31:0]    reg_activation_1_52;
wire signed[31:0]    reg_activation_1_53;
wire signed[31:0]    reg_activation_1_54;
wire signed[31:0]    reg_activation_1_55;
wire signed[31:0]    reg_activation_1_56;
wire signed[31:0]    reg_activation_1_57;
wire signed[31:0]    reg_activation_1_58;
wire signed[31:0]    reg_activation_1_59;
wire signed[31:0]    reg_activation_1_60;
wire signed[31:0]    reg_activation_1_61;
wire signed[31:0]    reg_activation_1_62;
wire signed[31:0]    reg_activation_1_63;
wire signed[31:0]    reg_activation_2_0;
wire signed[31:0]    reg_activation_2_1;
wire signed[31:0]    reg_activation_2_2;
wire signed[31:0]    reg_activation_2_3;
wire signed[31:0]    reg_activation_2_4;
wire signed[31:0]    reg_activation_2_5;
wire signed[31:0]    reg_activation_2_6;
wire signed[31:0]    reg_activation_2_7;
wire signed[31:0]    reg_activation_2_8;
wire signed[31:0]    reg_activation_2_9;
wire signed[31:0]    reg_activation_2_10;
wire signed[31:0]    reg_activation_2_11;
wire signed[31:0]    reg_activation_2_12;
wire signed[31:0]    reg_activation_2_13;
wire signed[31:0]    reg_activation_2_14;
wire signed[31:0]    reg_activation_2_15;
wire signed[31:0]    reg_activation_2_16;
wire signed[31:0]    reg_activation_2_17;
wire signed[31:0]    reg_activation_2_18;
wire signed[31:0]    reg_activation_2_19;
wire signed[31:0]    reg_activation_2_20;
wire signed[31:0]    reg_activation_2_21;
wire signed[31:0]    reg_activation_2_22;
wire signed[31:0]    reg_activation_2_23;
wire signed[31:0]    reg_activation_2_24;
wire signed[31:0]    reg_activation_2_25;
wire signed[31:0]    reg_activation_2_26;
wire signed[31:0]    reg_activation_2_27;
wire signed[31:0]    reg_activation_2_28;
wire signed[31:0]    reg_activation_2_29;
wire signed[31:0]    reg_activation_2_30;
wire signed[31:0]    reg_activation_2_31;
wire signed[31:0]    reg_activation_2_32;
wire signed[31:0]    reg_activation_2_33;
wire signed[31:0]    reg_activation_2_34;
wire signed[31:0]    reg_activation_2_35;
wire signed[31:0]    reg_activation_2_36;
wire signed[31:0]    reg_activation_2_37;
wire signed[31:0]    reg_activation_2_38;
wire signed[31:0]    reg_activation_2_39;
wire signed[31:0]    reg_activation_2_40;
wire signed[31:0]    reg_activation_2_41;
wire signed[31:0]    reg_activation_2_42;
wire signed[31:0]    reg_activation_2_43;
wire signed[31:0]    reg_activation_2_44;
wire signed[31:0]    reg_activation_2_45;
wire signed[31:0]    reg_activation_2_46;
wire signed[31:0]    reg_activation_2_47;
wire signed[31:0]    reg_activation_2_48;
wire signed[31:0]    reg_activation_2_49;
wire signed[31:0]    reg_activation_2_50;
wire signed[31:0]    reg_activation_2_51;
wire signed[31:0]    reg_activation_2_52;
wire signed[31:0]    reg_activation_2_53;
wire signed[31:0]    reg_activation_2_54;
wire signed[31:0]    reg_activation_2_55;
wire signed[31:0]    reg_activation_2_56;
wire signed[31:0]    reg_activation_2_57;
wire signed[31:0]    reg_activation_2_58;
wire signed[31:0]    reg_activation_2_59;
wire signed[31:0]    reg_activation_2_60;
wire signed[31:0]    reg_activation_2_61;
wire signed[31:0]    reg_activation_2_62;
wire signed[31:0]    reg_activation_2_63;
wire signed[31:0]    reg_activation_3_0;
wire signed[31:0]    reg_activation_3_1;
wire signed[31:0]    reg_activation_3_2;
wire signed[31:0]    reg_activation_3_3;
wire signed[31:0]    reg_activation_3_4;
wire signed[31:0]    reg_activation_3_5;
wire signed[31:0]    reg_activation_3_6;
wire signed[31:0]    reg_activation_3_7;
wire signed[31:0]    reg_activation_3_8;
wire signed[31:0]    reg_activation_3_9;
wire signed[31:0]    reg_activation_3_10;
wire signed[31:0]    reg_activation_3_11;
wire signed[31:0]    reg_activation_3_12;
wire signed[31:0]    reg_activation_3_13;
wire signed[31:0]    reg_activation_3_14;
wire signed[31:0]    reg_activation_3_15;
wire signed[31:0]    reg_activation_3_16;
wire signed[31:0]    reg_activation_3_17;
wire signed[31:0]    reg_activation_3_18;
wire signed[31:0]    reg_activation_3_19;
wire signed[31:0]    reg_activation_3_20;
wire signed[31:0]    reg_activation_3_21;
wire signed[31:0]    reg_activation_3_22;
wire signed[31:0]    reg_activation_3_23;
wire signed[31:0]    reg_activation_3_24;
wire signed[31:0]    reg_activation_3_25;
wire signed[31:0]    reg_activation_3_26;
wire signed[31:0]    reg_activation_3_27;
wire signed[31:0]    reg_activation_3_28;
wire signed[31:0]    reg_activation_3_29;
wire signed[31:0]    reg_activation_3_30;
wire signed[31:0]    reg_activation_3_31;
wire signed[31:0]    reg_activation_3_32;
wire signed[31:0]    reg_activation_3_33;
wire signed[31:0]    reg_activation_3_34;
wire signed[31:0]    reg_activation_3_35;
wire signed[31:0]    reg_activation_3_36;
wire signed[31:0]    reg_activation_3_37;
wire signed[31:0]    reg_activation_3_38;
wire signed[31:0]    reg_activation_3_39;
wire signed[31:0]    reg_activation_3_40;
wire signed[31:0]    reg_activation_3_41;
wire signed[31:0]    reg_activation_3_42;
wire signed[31:0]    reg_activation_3_43;
wire signed[31:0]    reg_activation_3_44;
wire signed[31:0]    reg_activation_3_45;
wire signed[31:0]    reg_activation_3_46;
wire signed[31:0]    reg_activation_3_47;
wire signed[31:0]    reg_activation_3_48;
wire signed[31:0]    reg_activation_3_49;
wire signed[31:0]    reg_activation_3_50;
wire signed[31:0]    reg_activation_3_51;
wire signed[31:0]    reg_activation_3_52;
wire signed[31:0]    reg_activation_3_53;
wire signed[31:0]    reg_activation_3_54;
wire signed[31:0]    reg_activation_3_55;
wire signed[31:0]    reg_activation_3_56;
wire signed[31:0]    reg_activation_3_57;
wire signed[31:0]    reg_activation_3_58;
wire signed[31:0]    reg_activation_3_59;
wire signed[31:0]    reg_activation_3_60;
wire signed[31:0]    reg_activation_3_61;
wire signed[31:0]    reg_activation_3_62;
wire signed[31:0]    reg_activation_3_63;
wire signed[31:0]    reg_activation_4_0;
wire signed[31:0]    reg_activation_4_1;
wire signed[31:0]    reg_activation_4_2;
wire signed[31:0]    reg_activation_4_3;
wire signed[31:0]    reg_activation_4_4;
wire signed[31:0]    reg_activation_4_5;
wire signed[31:0]    reg_activation_4_6;
wire signed[31:0]    reg_activation_4_7;
wire signed[31:0]    reg_activation_4_8;
wire signed[31:0]    reg_activation_4_9;
wire signed[31:0]    reg_activation_4_10;
wire signed[31:0]    reg_activation_4_11;
wire signed[31:0]    reg_activation_4_12;
wire signed[31:0]    reg_activation_4_13;
wire signed[31:0]    reg_activation_4_14;
wire signed[31:0]    reg_activation_4_15;
wire signed[31:0]    reg_activation_4_16;
wire signed[31:0]    reg_activation_4_17;
wire signed[31:0]    reg_activation_4_18;
wire signed[31:0]    reg_activation_4_19;
wire signed[31:0]    reg_activation_4_20;
wire signed[31:0]    reg_activation_4_21;
wire signed[31:0]    reg_activation_4_22;
wire signed[31:0]    reg_activation_4_23;
wire signed[31:0]    reg_activation_4_24;
wire signed[31:0]    reg_activation_4_25;
wire signed[31:0]    reg_activation_4_26;
wire signed[31:0]    reg_activation_4_27;
wire signed[31:0]    reg_activation_4_28;
wire signed[31:0]    reg_activation_4_29;
wire signed[31:0]    reg_activation_4_30;
wire signed[31:0]    reg_activation_4_31;
wire signed[31:0]    reg_activation_4_32;
wire signed[31:0]    reg_activation_4_33;
wire signed[31:0]    reg_activation_4_34;
wire signed[31:0]    reg_activation_4_35;
wire signed[31:0]    reg_activation_4_36;
wire signed[31:0]    reg_activation_4_37;
wire signed[31:0]    reg_activation_4_38;
wire signed[31:0]    reg_activation_4_39;
wire signed[31:0]    reg_activation_4_40;
wire signed[31:0]    reg_activation_4_41;
wire signed[31:0]    reg_activation_4_42;
wire signed[31:0]    reg_activation_4_43;
wire signed[31:0]    reg_activation_4_44;
wire signed[31:0]    reg_activation_4_45;
wire signed[31:0]    reg_activation_4_46;
wire signed[31:0]    reg_activation_4_47;
wire signed[31:0]    reg_activation_4_48;
wire signed[31:0]    reg_activation_4_49;
wire signed[31:0]    reg_activation_4_50;
wire signed[31:0]    reg_activation_4_51;
wire signed[31:0]    reg_activation_4_52;
wire signed[31:0]    reg_activation_4_53;
wire signed[31:0]    reg_activation_4_54;
wire signed[31:0]    reg_activation_4_55;
wire signed[31:0]    reg_activation_4_56;
wire signed[31:0]    reg_activation_4_57;
wire signed[31:0]    reg_activation_4_58;
wire signed[31:0]    reg_activation_4_59;
wire signed[31:0]    reg_activation_4_60;
wire signed[31:0]    reg_activation_4_61;
wire signed[31:0]    reg_activation_4_62;
wire signed[31:0]    reg_activation_4_63;
wire signed[31:0]    reg_activation_5_0;
wire signed[31:0]    reg_activation_5_1;
wire signed[31:0]    reg_activation_5_2;
wire signed[31:0]    reg_activation_5_3;
wire signed[31:0]    reg_activation_5_4;
wire signed[31:0]    reg_activation_5_5;
wire signed[31:0]    reg_activation_5_6;
wire signed[31:0]    reg_activation_5_7;
wire signed[31:0]    reg_activation_5_8;
wire signed[31:0]    reg_activation_5_9;
wire signed[31:0]    reg_activation_5_10;
wire signed[31:0]    reg_activation_5_11;
wire signed[31:0]    reg_activation_5_12;
wire signed[31:0]    reg_activation_5_13;
wire signed[31:0]    reg_activation_5_14;
wire signed[31:0]    reg_activation_5_15;
wire signed[31:0]    reg_activation_5_16;
wire signed[31:0]    reg_activation_5_17;
wire signed[31:0]    reg_activation_5_18;
wire signed[31:0]    reg_activation_5_19;
wire signed[31:0]    reg_activation_5_20;
wire signed[31:0]    reg_activation_5_21;
wire signed[31:0]    reg_activation_5_22;
wire signed[31:0]    reg_activation_5_23;
wire signed[31:0]    reg_activation_5_24;
wire signed[31:0]    reg_activation_5_25;
wire signed[31:0]    reg_activation_5_26;
wire signed[31:0]    reg_activation_5_27;
wire signed[31:0]    reg_activation_5_28;
wire signed[31:0]    reg_activation_5_29;
wire signed[31:0]    reg_activation_5_30;
wire signed[31:0]    reg_activation_5_31;
wire signed[31:0]    reg_activation_5_32;
wire signed[31:0]    reg_activation_5_33;
wire signed[31:0]    reg_activation_5_34;
wire signed[31:0]    reg_activation_5_35;
wire signed[31:0]    reg_activation_5_36;
wire signed[31:0]    reg_activation_5_37;
wire signed[31:0]    reg_activation_5_38;
wire signed[31:0]    reg_activation_5_39;
wire signed[31:0]    reg_activation_5_40;
wire signed[31:0]    reg_activation_5_41;
wire signed[31:0]    reg_activation_5_42;
wire signed[31:0]    reg_activation_5_43;
wire signed[31:0]    reg_activation_5_44;
wire signed[31:0]    reg_activation_5_45;
wire signed[31:0]    reg_activation_5_46;
wire signed[31:0]    reg_activation_5_47;
wire signed[31:0]    reg_activation_5_48;
wire signed[31:0]    reg_activation_5_49;
wire signed[31:0]    reg_activation_5_50;
wire signed[31:0]    reg_activation_5_51;
wire signed[31:0]    reg_activation_5_52;
wire signed[31:0]    reg_activation_5_53;
wire signed[31:0]    reg_activation_5_54;
wire signed[31:0]    reg_activation_5_55;
wire signed[31:0]    reg_activation_5_56;
wire signed[31:0]    reg_activation_5_57;
wire signed[31:0]    reg_activation_5_58;
wire signed[31:0]    reg_activation_5_59;
wire signed[31:0]    reg_activation_5_60;
wire signed[31:0]    reg_activation_5_61;
wire signed[31:0]    reg_activation_5_62;
wire signed[31:0]    reg_activation_5_63;
wire signed[31:0]    reg_activation_6_0;
wire signed[31:0]    reg_activation_6_1;
wire signed[31:0]    reg_activation_6_2;
wire signed[31:0]    reg_activation_6_3;
wire signed[31:0]    reg_activation_6_4;
wire signed[31:0]    reg_activation_6_5;
wire signed[31:0]    reg_activation_6_6;
wire signed[31:0]    reg_activation_6_7;
wire signed[31:0]    reg_activation_6_8;
wire signed[31:0]    reg_activation_6_9;
wire signed[31:0]    reg_activation_6_10;
wire signed[31:0]    reg_activation_6_11;
wire signed[31:0]    reg_activation_6_12;
wire signed[31:0]    reg_activation_6_13;
wire signed[31:0]    reg_activation_6_14;
wire signed[31:0]    reg_activation_6_15;
wire signed[31:0]    reg_activation_6_16;
wire signed[31:0]    reg_activation_6_17;
wire signed[31:0]    reg_activation_6_18;
wire signed[31:0]    reg_activation_6_19;
wire signed[31:0]    reg_activation_6_20;
wire signed[31:0]    reg_activation_6_21;
wire signed[31:0]    reg_activation_6_22;
wire signed[31:0]    reg_activation_6_23;
wire signed[31:0]    reg_activation_6_24;
wire signed[31:0]    reg_activation_6_25;
wire signed[31:0]    reg_activation_6_26;
wire signed[31:0]    reg_activation_6_27;
wire signed[31:0]    reg_activation_6_28;
wire signed[31:0]    reg_activation_6_29;
wire signed[31:0]    reg_activation_6_30;
wire signed[31:0]    reg_activation_6_31;
wire signed[31:0]    reg_activation_6_32;
wire signed[31:0]    reg_activation_6_33;
wire signed[31:0]    reg_activation_6_34;
wire signed[31:0]    reg_activation_6_35;
wire signed[31:0]    reg_activation_6_36;
wire signed[31:0]    reg_activation_6_37;
wire signed[31:0]    reg_activation_6_38;
wire signed[31:0]    reg_activation_6_39;
wire signed[31:0]    reg_activation_6_40;
wire signed[31:0]    reg_activation_6_41;
wire signed[31:0]    reg_activation_6_42;
wire signed[31:0]    reg_activation_6_43;
wire signed[31:0]    reg_activation_6_44;
wire signed[31:0]    reg_activation_6_45;
wire signed[31:0]    reg_activation_6_46;
wire signed[31:0]    reg_activation_6_47;
wire signed[31:0]    reg_activation_6_48;
wire signed[31:0]    reg_activation_6_49;
wire signed[31:0]    reg_activation_6_50;
wire signed[31:0]    reg_activation_6_51;
wire signed[31:0]    reg_activation_6_52;
wire signed[31:0]    reg_activation_6_53;
wire signed[31:0]    reg_activation_6_54;
wire signed[31:0]    reg_activation_6_55;
wire signed[31:0]    reg_activation_6_56;
wire signed[31:0]    reg_activation_6_57;
wire signed[31:0]    reg_activation_6_58;
wire signed[31:0]    reg_activation_6_59;
wire signed[31:0]    reg_activation_6_60;
wire signed[31:0]    reg_activation_6_61;
wire signed[31:0]    reg_activation_6_62;
wire signed[31:0]    reg_activation_6_63;
wire signed[31:0]    reg_activation_7_0;
wire signed[31:0]    reg_activation_7_1;
wire signed[31:0]    reg_activation_7_2;
wire signed[31:0]    reg_activation_7_3;
wire signed[31:0]    reg_activation_7_4;
wire signed[31:0]    reg_activation_7_5;
wire signed[31:0]    reg_activation_7_6;
wire signed[31:0]    reg_activation_7_7;
wire signed[31:0]    reg_activation_7_8;
wire signed[31:0]    reg_activation_7_9;
wire signed[31:0]    reg_activation_7_10;
wire signed[31:0]    reg_activation_7_11;
wire signed[31:0]    reg_activation_7_12;
wire signed[31:0]    reg_activation_7_13;
wire signed[31:0]    reg_activation_7_14;
wire signed[31:0]    reg_activation_7_15;
wire signed[31:0]    reg_activation_7_16;
wire signed[31:0]    reg_activation_7_17;
wire signed[31:0]    reg_activation_7_18;
wire signed[31:0]    reg_activation_7_19;
wire signed[31:0]    reg_activation_7_20;
wire signed[31:0]    reg_activation_7_21;
wire signed[31:0]    reg_activation_7_22;
wire signed[31:0]    reg_activation_7_23;
wire signed[31:0]    reg_activation_7_24;
wire signed[31:0]    reg_activation_7_25;
wire signed[31:0]    reg_activation_7_26;
wire signed[31:0]    reg_activation_7_27;
wire signed[31:0]    reg_activation_7_28;
wire signed[31:0]    reg_activation_7_29;
wire signed[31:0]    reg_activation_7_30;
wire signed[31:0]    reg_activation_7_31;
wire signed[31:0]    reg_activation_7_32;
wire signed[31:0]    reg_activation_7_33;
wire signed[31:0]    reg_activation_7_34;
wire signed[31:0]    reg_activation_7_35;
wire signed[31:0]    reg_activation_7_36;
wire signed[31:0]    reg_activation_7_37;
wire signed[31:0]    reg_activation_7_38;
wire signed[31:0]    reg_activation_7_39;
wire signed[31:0]    reg_activation_7_40;
wire signed[31:0]    reg_activation_7_41;
wire signed[31:0]    reg_activation_7_42;
wire signed[31:0]    reg_activation_7_43;
wire signed[31:0]    reg_activation_7_44;
wire signed[31:0]    reg_activation_7_45;
wire signed[31:0]    reg_activation_7_46;
wire signed[31:0]    reg_activation_7_47;
wire signed[31:0]    reg_activation_7_48;
wire signed[31:0]    reg_activation_7_49;
wire signed[31:0]    reg_activation_7_50;
wire signed[31:0]    reg_activation_7_51;
wire signed[31:0]    reg_activation_7_52;
wire signed[31:0]    reg_activation_7_53;
wire signed[31:0]    reg_activation_7_54;
wire signed[31:0]    reg_activation_7_55;
wire signed[31:0]    reg_activation_7_56;
wire signed[31:0]    reg_activation_7_57;
wire signed[31:0]    reg_activation_7_58;
wire signed[31:0]    reg_activation_7_59;
wire signed[31:0]    reg_activation_7_60;
wire signed[31:0]    reg_activation_7_61;
wire signed[31:0]    reg_activation_7_62;
wire signed[31:0]    reg_activation_7_63;
wire signed[31:0]    reg_activation_8_0;
wire signed[31:0]    reg_activation_8_1;
wire signed[31:0]    reg_activation_8_2;
wire signed[31:0]    reg_activation_8_3;
wire signed[31:0]    reg_activation_8_4;
wire signed[31:0]    reg_activation_8_5;
wire signed[31:0]    reg_activation_8_6;
wire signed[31:0]    reg_activation_8_7;
wire signed[31:0]    reg_activation_8_8;
wire signed[31:0]    reg_activation_8_9;
wire signed[31:0]    reg_activation_8_10;
wire signed[31:0]    reg_activation_8_11;
wire signed[31:0]    reg_activation_8_12;
wire signed[31:0]    reg_activation_8_13;
wire signed[31:0]    reg_activation_8_14;
wire signed[31:0]    reg_activation_8_15;
wire signed[31:0]    reg_activation_8_16;
wire signed[31:0]    reg_activation_8_17;
wire signed[31:0]    reg_activation_8_18;
wire signed[31:0]    reg_activation_8_19;
wire signed[31:0]    reg_activation_8_20;
wire signed[31:0]    reg_activation_8_21;
wire signed[31:0]    reg_activation_8_22;
wire signed[31:0]    reg_activation_8_23;
wire signed[31:0]    reg_activation_8_24;
wire signed[31:0]    reg_activation_8_25;
wire signed[31:0]    reg_activation_8_26;
wire signed[31:0]    reg_activation_8_27;
wire signed[31:0]    reg_activation_8_28;
wire signed[31:0]    reg_activation_8_29;
wire signed[31:0]    reg_activation_8_30;
wire signed[31:0]    reg_activation_8_31;
wire signed[31:0]    reg_activation_8_32;
wire signed[31:0]    reg_activation_8_33;
wire signed[31:0]    reg_activation_8_34;
wire signed[31:0]    reg_activation_8_35;
wire signed[31:0]    reg_activation_8_36;
wire signed[31:0]    reg_activation_8_37;
wire signed[31:0]    reg_activation_8_38;
wire signed[31:0]    reg_activation_8_39;
wire signed[31:0]    reg_activation_8_40;
wire signed[31:0]    reg_activation_8_41;
wire signed[31:0]    reg_activation_8_42;
wire signed[31:0]    reg_activation_8_43;
wire signed[31:0]    reg_activation_8_44;
wire signed[31:0]    reg_activation_8_45;
wire signed[31:0]    reg_activation_8_46;
wire signed[31:0]    reg_activation_8_47;
wire signed[31:0]    reg_activation_8_48;
wire signed[31:0]    reg_activation_8_49;
wire signed[31:0]    reg_activation_8_50;
wire signed[31:0]    reg_activation_8_51;
wire signed[31:0]    reg_activation_8_52;
wire signed[31:0]    reg_activation_8_53;
wire signed[31:0]    reg_activation_8_54;
wire signed[31:0]    reg_activation_8_55;
wire signed[31:0]    reg_activation_8_56;
wire signed[31:0]    reg_activation_8_57;
wire signed[31:0]    reg_activation_8_58;
wire signed[31:0]    reg_activation_8_59;
wire signed[31:0]    reg_activation_8_60;
wire signed[31:0]    reg_activation_8_61;
wire signed[31:0]    reg_activation_8_62;
wire signed[31:0]    reg_activation_8_63;
wire signed[31:0]    reg_activation_9_0;
wire signed[31:0]    reg_activation_9_1;
wire signed[31:0]    reg_activation_9_2;
wire signed[31:0]    reg_activation_9_3;
wire signed[31:0]    reg_activation_9_4;
wire signed[31:0]    reg_activation_9_5;
wire signed[31:0]    reg_activation_9_6;
wire signed[31:0]    reg_activation_9_7;
wire signed[31:0]    reg_activation_9_8;
wire signed[31:0]    reg_activation_9_9;
wire signed[31:0]    reg_activation_9_10;
wire signed[31:0]    reg_activation_9_11;
wire signed[31:0]    reg_activation_9_12;
wire signed[31:0]    reg_activation_9_13;
wire signed[31:0]    reg_activation_9_14;
wire signed[31:0]    reg_activation_9_15;
wire signed[31:0]    reg_activation_9_16;
wire signed[31:0]    reg_activation_9_17;
wire signed[31:0]    reg_activation_9_18;
wire signed[31:0]    reg_activation_9_19;
wire signed[31:0]    reg_activation_9_20;
wire signed[31:0]    reg_activation_9_21;
wire signed[31:0]    reg_activation_9_22;
wire signed[31:0]    reg_activation_9_23;
wire signed[31:0]    reg_activation_9_24;
wire signed[31:0]    reg_activation_9_25;
wire signed[31:0]    reg_activation_9_26;
wire signed[31:0]    reg_activation_9_27;
wire signed[31:0]    reg_activation_9_28;
wire signed[31:0]    reg_activation_9_29;
wire signed[31:0]    reg_activation_9_30;
wire signed[31:0]    reg_activation_9_31;
wire signed[31:0]    reg_activation_9_32;
wire signed[31:0]    reg_activation_9_33;
wire signed[31:0]    reg_activation_9_34;
wire signed[31:0]    reg_activation_9_35;
wire signed[31:0]    reg_activation_9_36;
wire signed[31:0]    reg_activation_9_37;
wire signed[31:0]    reg_activation_9_38;
wire signed[31:0]    reg_activation_9_39;
wire signed[31:0]    reg_activation_9_40;
wire signed[31:0]    reg_activation_9_41;
wire signed[31:0]    reg_activation_9_42;
wire signed[31:0]    reg_activation_9_43;
wire signed[31:0]    reg_activation_9_44;
wire signed[31:0]    reg_activation_9_45;
wire signed[31:0]    reg_activation_9_46;
wire signed[31:0]    reg_activation_9_47;
wire signed[31:0]    reg_activation_9_48;
wire signed[31:0]    reg_activation_9_49;
wire signed[31:0]    reg_activation_9_50;
wire signed[31:0]    reg_activation_9_51;
wire signed[31:0]    reg_activation_9_52;
wire signed[31:0]    reg_activation_9_53;
wire signed[31:0]    reg_activation_9_54;
wire signed[31:0]    reg_activation_9_55;
wire signed[31:0]    reg_activation_9_56;
wire signed[31:0]    reg_activation_9_57;
wire signed[31:0]    reg_activation_9_58;
wire signed[31:0]    reg_activation_9_59;
wire signed[31:0]    reg_activation_9_60;
wire signed[31:0]    reg_activation_9_61;
wire signed[31:0]    reg_activation_9_62;
wire signed[31:0]    reg_activation_9_63;
wire signed[31:0]    reg_activation_10_0;
wire signed[31:0]    reg_activation_10_1;
wire signed[31:0]    reg_activation_10_2;
wire signed[31:0]    reg_activation_10_3;
wire signed[31:0]    reg_activation_10_4;
wire signed[31:0]    reg_activation_10_5;
wire signed[31:0]    reg_activation_10_6;
wire signed[31:0]    reg_activation_10_7;
wire signed[31:0]    reg_activation_10_8;
wire signed[31:0]    reg_activation_10_9;
wire signed[31:0]    reg_activation_10_10;
wire signed[31:0]    reg_activation_10_11;
wire signed[31:0]    reg_activation_10_12;
wire signed[31:0]    reg_activation_10_13;
wire signed[31:0]    reg_activation_10_14;
wire signed[31:0]    reg_activation_10_15;
wire signed[31:0]    reg_activation_10_16;
wire signed[31:0]    reg_activation_10_17;
wire signed[31:0]    reg_activation_10_18;
wire signed[31:0]    reg_activation_10_19;
wire signed[31:0]    reg_activation_10_20;
wire signed[31:0]    reg_activation_10_21;
wire signed[31:0]    reg_activation_10_22;
wire signed[31:0]    reg_activation_10_23;
wire signed[31:0]    reg_activation_10_24;
wire signed[31:0]    reg_activation_10_25;
wire signed[31:0]    reg_activation_10_26;
wire signed[31:0]    reg_activation_10_27;
wire signed[31:0]    reg_activation_10_28;
wire signed[31:0]    reg_activation_10_29;
wire signed[31:0]    reg_activation_10_30;
wire signed[31:0]    reg_activation_10_31;
wire signed[31:0]    reg_activation_10_32;
wire signed[31:0]    reg_activation_10_33;
wire signed[31:0]    reg_activation_10_34;
wire signed[31:0]    reg_activation_10_35;
wire signed[31:0]    reg_activation_10_36;
wire signed[31:0]    reg_activation_10_37;
wire signed[31:0]    reg_activation_10_38;
wire signed[31:0]    reg_activation_10_39;
wire signed[31:0]    reg_activation_10_40;
wire signed[31:0]    reg_activation_10_41;
wire signed[31:0]    reg_activation_10_42;
wire signed[31:0]    reg_activation_10_43;
wire signed[31:0]    reg_activation_10_44;
wire signed[31:0]    reg_activation_10_45;
wire signed[31:0]    reg_activation_10_46;
wire signed[31:0]    reg_activation_10_47;
wire signed[31:0]    reg_activation_10_48;
wire signed[31:0]    reg_activation_10_49;
wire signed[31:0]    reg_activation_10_50;
wire signed[31:0]    reg_activation_10_51;
wire signed[31:0]    reg_activation_10_52;
wire signed[31:0]    reg_activation_10_53;
wire signed[31:0]    reg_activation_10_54;
wire signed[31:0]    reg_activation_10_55;
wire signed[31:0]    reg_activation_10_56;
wire signed[31:0]    reg_activation_10_57;
wire signed[31:0]    reg_activation_10_58;
wire signed[31:0]    reg_activation_10_59;
wire signed[31:0]    reg_activation_10_60;
wire signed[31:0]    reg_activation_10_61;
wire signed[31:0]    reg_activation_10_62;
wire signed[31:0]    reg_activation_10_63;
wire signed[31:0]    reg_activation_11_0;
wire signed[31:0]    reg_activation_11_1;
wire signed[31:0]    reg_activation_11_2;
wire signed[31:0]    reg_activation_11_3;
wire signed[31:0]    reg_activation_11_4;
wire signed[31:0]    reg_activation_11_5;
wire signed[31:0]    reg_activation_11_6;
wire signed[31:0]    reg_activation_11_7;
wire signed[31:0]    reg_activation_11_8;
wire signed[31:0]    reg_activation_11_9;
wire signed[31:0]    reg_activation_11_10;
wire signed[31:0]    reg_activation_11_11;
wire signed[31:0]    reg_activation_11_12;
wire signed[31:0]    reg_activation_11_13;
wire signed[31:0]    reg_activation_11_14;
wire signed[31:0]    reg_activation_11_15;
wire signed[31:0]    reg_activation_11_16;
wire signed[31:0]    reg_activation_11_17;
wire signed[31:0]    reg_activation_11_18;
wire signed[31:0]    reg_activation_11_19;
wire signed[31:0]    reg_activation_11_20;
wire signed[31:0]    reg_activation_11_21;
wire signed[31:0]    reg_activation_11_22;
wire signed[31:0]    reg_activation_11_23;
wire signed[31:0]    reg_activation_11_24;
wire signed[31:0]    reg_activation_11_25;
wire signed[31:0]    reg_activation_11_26;
wire signed[31:0]    reg_activation_11_27;
wire signed[31:0]    reg_activation_11_28;
wire signed[31:0]    reg_activation_11_29;
wire signed[31:0]    reg_activation_11_30;
wire signed[31:0]    reg_activation_11_31;
wire signed[31:0]    reg_activation_11_32;
wire signed[31:0]    reg_activation_11_33;
wire signed[31:0]    reg_activation_11_34;
wire signed[31:0]    reg_activation_11_35;
wire signed[31:0]    reg_activation_11_36;
wire signed[31:0]    reg_activation_11_37;
wire signed[31:0]    reg_activation_11_38;
wire signed[31:0]    reg_activation_11_39;
wire signed[31:0]    reg_activation_11_40;
wire signed[31:0]    reg_activation_11_41;
wire signed[31:0]    reg_activation_11_42;
wire signed[31:0]    reg_activation_11_43;
wire signed[31:0]    reg_activation_11_44;
wire signed[31:0]    reg_activation_11_45;
wire signed[31:0]    reg_activation_11_46;
wire signed[31:0]    reg_activation_11_47;
wire signed[31:0]    reg_activation_11_48;
wire signed[31:0]    reg_activation_11_49;
wire signed[31:0]    reg_activation_11_50;
wire signed[31:0]    reg_activation_11_51;
wire signed[31:0]    reg_activation_11_52;
wire signed[31:0]    reg_activation_11_53;
wire signed[31:0]    reg_activation_11_54;
wire signed[31:0]    reg_activation_11_55;
wire signed[31:0]    reg_activation_11_56;
wire signed[31:0]    reg_activation_11_57;
wire signed[31:0]    reg_activation_11_58;
wire signed[31:0]    reg_activation_11_59;
wire signed[31:0]    reg_activation_11_60;
wire signed[31:0]    reg_activation_11_61;
wire signed[31:0]    reg_activation_11_62;
wire signed[31:0]    reg_activation_11_63;
wire signed[31:0]    reg_activation_12_0;
wire signed[31:0]    reg_activation_12_1;
wire signed[31:0]    reg_activation_12_2;
wire signed[31:0]    reg_activation_12_3;
wire signed[31:0]    reg_activation_12_4;
wire signed[31:0]    reg_activation_12_5;
wire signed[31:0]    reg_activation_12_6;
wire signed[31:0]    reg_activation_12_7;
wire signed[31:0]    reg_activation_12_8;
wire signed[31:0]    reg_activation_12_9;
wire signed[31:0]    reg_activation_12_10;
wire signed[31:0]    reg_activation_12_11;
wire signed[31:0]    reg_activation_12_12;
wire signed[31:0]    reg_activation_12_13;
wire signed[31:0]    reg_activation_12_14;
wire signed[31:0]    reg_activation_12_15;
wire signed[31:0]    reg_activation_12_16;
wire signed[31:0]    reg_activation_12_17;
wire signed[31:0]    reg_activation_12_18;
wire signed[31:0]    reg_activation_12_19;
wire signed[31:0]    reg_activation_12_20;
wire signed[31:0]    reg_activation_12_21;
wire signed[31:0]    reg_activation_12_22;
wire signed[31:0]    reg_activation_12_23;
wire signed[31:0]    reg_activation_12_24;
wire signed[31:0]    reg_activation_12_25;
wire signed[31:0]    reg_activation_12_26;
wire signed[31:0]    reg_activation_12_27;
wire signed[31:0]    reg_activation_12_28;
wire signed[31:0]    reg_activation_12_29;
wire signed[31:0]    reg_activation_12_30;
wire signed[31:0]    reg_activation_12_31;
wire signed[31:0]    reg_activation_12_32;
wire signed[31:0]    reg_activation_12_33;
wire signed[31:0]    reg_activation_12_34;
wire signed[31:0]    reg_activation_12_35;
wire signed[31:0]    reg_activation_12_36;
wire signed[31:0]    reg_activation_12_37;
wire signed[31:0]    reg_activation_12_38;
wire signed[31:0]    reg_activation_12_39;
wire signed[31:0]    reg_activation_12_40;
wire signed[31:0]    reg_activation_12_41;
wire signed[31:0]    reg_activation_12_42;
wire signed[31:0]    reg_activation_12_43;
wire signed[31:0]    reg_activation_12_44;
wire signed[31:0]    reg_activation_12_45;
wire signed[31:0]    reg_activation_12_46;
wire signed[31:0]    reg_activation_12_47;
wire signed[31:0]    reg_activation_12_48;
wire signed[31:0]    reg_activation_12_49;
wire signed[31:0]    reg_activation_12_50;
wire signed[31:0]    reg_activation_12_51;
wire signed[31:0]    reg_activation_12_52;
wire signed[31:0]    reg_activation_12_53;
wire signed[31:0]    reg_activation_12_54;
wire signed[31:0]    reg_activation_12_55;
wire signed[31:0]    reg_activation_12_56;
wire signed[31:0]    reg_activation_12_57;
wire signed[31:0]    reg_activation_12_58;
wire signed[31:0]    reg_activation_12_59;
wire signed[31:0]    reg_activation_12_60;
wire signed[31:0]    reg_activation_12_61;
wire signed[31:0]    reg_activation_12_62;
wire signed[31:0]    reg_activation_12_63;
wire signed[31:0]    reg_activation_13_0;
wire signed[31:0]    reg_activation_13_1;
wire signed[31:0]    reg_activation_13_2;
wire signed[31:0]    reg_activation_13_3;
wire signed[31:0]    reg_activation_13_4;
wire signed[31:0]    reg_activation_13_5;
wire signed[31:0]    reg_activation_13_6;
wire signed[31:0]    reg_activation_13_7;
wire signed[31:0]    reg_activation_13_8;
wire signed[31:0]    reg_activation_13_9;
wire signed[31:0]    reg_activation_13_10;
wire signed[31:0]    reg_activation_13_11;
wire signed[31:0]    reg_activation_13_12;
wire signed[31:0]    reg_activation_13_13;
wire signed[31:0]    reg_activation_13_14;
wire signed[31:0]    reg_activation_13_15;
wire signed[31:0]    reg_activation_13_16;
wire signed[31:0]    reg_activation_13_17;
wire signed[31:0]    reg_activation_13_18;
wire signed[31:0]    reg_activation_13_19;
wire signed[31:0]    reg_activation_13_20;
wire signed[31:0]    reg_activation_13_21;
wire signed[31:0]    reg_activation_13_22;
wire signed[31:0]    reg_activation_13_23;
wire signed[31:0]    reg_activation_13_24;
wire signed[31:0]    reg_activation_13_25;
wire signed[31:0]    reg_activation_13_26;
wire signed[31:0]    reg_activation_13_27;
wire signed[31:0]    reg_activation_13_28;
wire signed[31:0]    reg_activation_13_29;
wire signed[31:0]    reg_activation_13_30;
wire signed[31:0]    reg_activation_13_31;
wire signed[31:0]    reg_activation_13_32;
wire signed[31:0]    reg_activation_13_33;
wire signed[31:0]    reg_activation_13_34;
wire signed[31:0]    reg_activation_13_35;
wire signed[31:0]    reg_activation_13_36;
wire signed[31:0]    reg_activation_13_37;
wire signed[31:0]    reg_activation_13_38;
wire signed[31:0]    reg_activation_13_39;
wire signed[31:0]    reg_activation_13_40;
wire signed[31:0]    reg_activation_13_41;
wire signed[31:0]    reg_activation_13_42;
wire signed[31:0]    reg_activation_13_43;
wire signed[31:0]    reg_activation_13_44;
wire signed[31:0]    reg_activation_13_45;
wire signed[31:0]    reg_activation_13_46;
wire signed[31:0]    reg_activation_13_47;
wire signed[31:0]    reg_activation_13_48;
wire signed[31:0]    reg_activation_13_49;
wire signed[31:0]    reg_activation_13_50;
wire signed[31:0]    reg_activation_13_51;
wire signed[31:0]    reg_activation_13_52;
wire signed[31:0]    reg_activation_13_53;
wire signed[31:0]    reg_activation_13_54;
wire signed[31:0]    reg_activation_13_55;
wire signed[31:0]    reg_activation_13_56;
wire signed[31:0]    reg_activation_13_57;
wire signed[31:0]    reg_activation_13_58;
wire signed[31:0]    reg_activation_13_59;
wire signed[31:0]    reg_activation_13_60;
wire signed[31:0]    reg_activation_13_61;
wire signed[31:0]    reg_activation_13_62;
wire signed[31:0]    reg_activation_13_63;
wire signed[31:0]    reg_activation_14_0;
wire signed[31:0]    reg_activation_14_1;
wire signed[31:0]    reg_activation_14_2;
wire signed[31:0]    reg_activation_14_3;
wire signed[31:0]    reg_activation_14_4;
wire signed[31:0]    reg_activation_14_5;
wire signed[31:0]    reg_activation_14_6;
wire signed[31:0]    reg_activation_14_7;
wire signed[31:0]    reg_activation_14_8;
wire signed[31:0]    reg_activation_14_9;
wire signed[31:0]    reg_activation_14_10;
wire signed[31:0]    reg_activation_14_11;
wire signed[31:0]    reg_activation_14_12;
wire signed[31:0]    reg_activation_14_13;
wire signed[31:0]    reg_activation_14_14;
wire signed[31:0]    reg_activation_14_15;
wire signed[31:0]    reg_activation_14_16;
wire signed[31:0]    reg_activation_14_17;
wire signed[31:0]    reg_activation_14_18;
wire signed[31:0]    reg_activation_14_19;
wire signed[31:0]    reg_activation_14_20;
wire signed[31:0]    reg_activation_14_21;
wire signed[31:0]    reg_activation_14_22;
wire signed[31:0]    reg_activation_14_23;
wire signed[31:0]    reg_activation_14_24;
wire signed[31:0]    reg_activation_14_25;
wire signed[31:0]    reg_activation_14_26;
wire signed[31:0]    reg_activation_14_27;
wire signed[31:0]    reg_activation_14_28;
wire signed[31:0]    reg_activation_14_29;
wire signed[31:0]    reg_activation_14_30;
wire signed[31:0]    reg_activation_14_31;
wire signed[31:0]    reg_activation_14_32;
wire signed[31:0]    reg_activation_14_33;
wire signed[31:0]    reg_activation_14_34;
wire signed[31:0]    reg_activation_14_35;
wire signed[31:0]    reg_activation_14_36;
wire signed[31:0]    reg_activation_14_37;
wire signed[31:0]    reg_activation_14_38;
wire signed[31:0]    reg_activation_14_39;
wire signed[31:0]    reg_activation_14_40;
wire signed[31:0]    reg_activation_14_41;
wire signed[31:0]    reg_activation_14_42;
wire signed[31:0]    reg_activation_14_43;
wire signed[31:0]    reg_activation_14_44;
wire signed[31:0]    reg_activation_14_45;
wire signed[31:0]    reg_activation_14_46;
wire signed[31:0]    reg_activation_14_47;
wire signed[31:0]    reg_activation_14_48;
wire signed[31:0]    reg_activation_14_49;
wire signed[31:0]    reg_activation_14_50;
wire signed[31:0]    reg_activation_14_51;
wire signed[31:0]    reg_activation_14_52;
wire signed[31:0]    reg_activation_14_53;
wire signed[31:0]    reg_activation_14_54;
wire signed[31:0]    reg_activation_14_55;
wire signed[31:0]    reg_activation_14_56;
wire signed[31:0]    reg_activation_14_57;
wire signed[31:0]    reg_activation_14_58;
wire signed[31:0]    reg_activation_14_59;
wire signed[31:0]    reg_activation_14_60;
wire signed[31:0]    reg_activation_14_61;
wire signed[31:0]    reg_activation_14_62;
wire signed[31:0]    reg_activation_14_63;
wire signed[31:0]    reg_activation_15_0;
wire signed[31:0]    reg_activation_15_1;
wire signed[31:0]    reg_activation_15_2;
wire signed[31:0]    reg_activation_15_3;
wire signed[31:0]    reg_activation_15_4;
wire signed[31:0]    reg_activation_15_5;
wire signed[31:0]    reg_activation_15_6;
wire signed[31:0]    reg_activation_15_7;
wire signed[31:0]    reg_activation_15_8;
wire signed[31:0]    reg_activation_15_9;
wire signed[31:0]    reg_activation_15_10;
wire signed[31:0]    reg_activation_15_11;
wire signed[31:0]    reg_activation_15_12;
wire signed[31:0]    reg_activation_15_13;
wire signed[31:0]    reg_activation_15_14;
wire signed[31:0]    reg_activation_15_15;
wire signed[31:0]    reg_activation_15_16;
wire signed[31:0]    reg_activation_15_17;
wire signed[31:0]    reg_activation_15_18;
wire signed[31:0]    reg_activation_15_19;
wire signed[31:0]    reg_activation_15_20;
wire signed[31:0]    reg_activation_15_21;
wire signed[31:0]    reg_activation_15_22;
wire signed[31:0]    reg_activation_15_23;
wire signed[31:0]    reg_activation_15_24;
wire signed[31:0]    reg_activation_15_25;
wire signed[31:0]    reg_activation_15_26;
wire signed[31:0]    reg_activation_15_27;
wire signed[31:0]    reg_activation_15_28;
wire signed[31:0]    reg_activation_15_29;
wire signed[31:0]    reg_activation_15_30;
wire signed[31:0]    reg_activation_15_31;
wire signed[31:0]    reg_activation_15_32;
wire signed[31:0]    reg_activation_15_33;
wire signed[31:0]    reg_activation_15_34;
wire signed[31:0]    reg_activation_15_35;
wire signed[31:0]    reg_activation_15_36;
wire signed[31:0]    reg_activation_15_37;
wire signed[31:0]    reg_activation_15_38;
wire signed[31:0]    reg_activation_15_39;
wire signed[31:0]    reg_activation_15_40;
wire signed[31:0]    reg_activation_15_41;
wire signed[31:0]    reg_activation_15_42;
wire signed[31:0]    reg_activation_15_43;
wire signed[31:0]    reg_activation_15_44;
wire signed[31:0]    reg_activation_15_45;
wire signed[31:0]    reg_activation_15_46;
wire signed[31:0]    reg_activation_15_47;
wire signed[31:0]    reg_activation_15_48;
wire signed[31:0]    reg_activation_15_49;
wire signed[31:0]    reg_activation_15_50;
wire signed[31:0]    reg_activation_15_51;
wire signed[31:0]    reg_activation_15_52;
wire signed[31:0]    reg_activation_15_53;
wire signed[31:0]    reg_activation_15_54;
wire signed[31:0]    reg_activation_15_55;
wire signed[31:0]    reg_activation_15_56;
wire signed[31:0]    reg_activation_15_57;
wire signed[31:0]    reg_activation_15_58;
wire signed[31:0]    reg_activation_15_59;
wire signed[31:0]    reg_activation_15_60;
wire signed[31:0]    reg_activation_15_61;
wire signed[31:0]    reg_activation_15_62;
wire signed[31:0]    reg_activation_15_63;
wire signed[31:0]    reg_activation_16_0;
wire signed[31:0]    reg_activation_16_1;
wire signed[31:0]    reg_activation_16_2;
wire signed[31:0]    reg_activation_16_3;
wire signed[31:0]    reg_activation_16_4;
wire signed[31:0]    reg_activation_16_5;
wire signed[31:0]    reg_activation_16_6;
wire signed[31:0]    reg_activation_16_7;
wire signed[31:0]    reg_activation_16_8;
wire signed[31:0]    reg_activation_16_9;
wire signed[31:0]    reg_activation_16_10;
wire signed[31:0]    reg_activation_16_11;
wire signed[31:0]    reg_activation_16_12;
wire signed[31:0]    reg_activation_16_13;
wire signed[31:0]    reg_activation_16_14;
wire signed[31:0]    reg_activation_16_15;
wire signed[31:0]    reg_activation_16_16;
wire signed[31:0]    reg_activation_16_17;
wire signed[31:0]    reg_activation_16_18;
wire signed[31:0]    reg_activation_16_19;
wire signed[31:0]    reg_activation_16_20;
wire signed[31:0]    reg_activation_16_21;
wire signed[31:0]    reg_activation_16_22;
wire signed[31:0]    reg_activation_16_23;
wire signed[31:0]    reg_activation_16_24;
wire signed[31:0]    reg_activation_16_25;
wire signed[31:0]    reg_activation_16_26;
wire signed[31:0]    reg_activation_16_27;
wire signed[31:0]    reg_activation_16_28;
wire signed[31:0]    reg_activation_16_29;
wire signed[31:0]    reg_activation_16_30;
wire signed[31:0]    reg_activation_16_31;
wire signed[31:0]    reg_activation_16_32;
wire signed[31:0]    reg_activation_16_33;
wire signed[31:0]    reg_activation_16_34;
wire signed[31:0]    reg_activation_16_35;
wire signed[31:0]    reg_activation_16_36;
wire signed[31:0]    reg_activation_16_37;
wire signed[31:0]    reg_activation_16_38;
wire signed[31:0]    reg_activation_16_39;
wire signed[31:0]    reg_activation_16_40;
wire signed[31:0]    reg_activation_16_41;
wire signed[31:0]    reg_activation_16_42;
wire signed[31:0]    reg_activation_16_43;
wire signed[31:0]    reg_activation_16_44;
wire signed[31:0]    reg_activation_16_45;
wire signed[31:0]    reg_activation_16_46;
wire signed[31:0]    reg_activation_16_47;
wire signed[31:0]    reg_activation_16_48;
wire signed[31:0]    reg_activation_16_49;
wire signed[31:0]    reg_activation_16_50;
wire signed[31:0]    reg_activation_16_51;
wire signed[31:0]    reg_activation_16_52;
wire signed[31:0]    reg_activation_16_53;
wire signed[31:0]    reg_activation_16_54;
wire signed[31:0]    reg_activation_16_55;
wire signed[31:0]    reg_activation_16_56;
wire signed[31:0]    reg_activation_16_57;
wire signed[31:0]    reg_activation_16_58;
wire signed[31:0]    reg_activation_16_59;
wire signed[31:0]    reg_activation_16_60;
wire signed[31:0]    reg_activation_16_61;
wire signed[31:0]    reg_activation_16_62;
wire signed[31:0]    reg_activation_16_63;
wire signed[31:0]    reg_activation_17_0;
wire signed[31:0]    reg_activation_17_1;
wire signed[31:0]    reg_activation_17_2;
wire signed[31:0]    reg_activation_17_3;
wire signed[31:0]    reg_activation_17_4;
wire signed[31:0]    reg_activation_17_5;
wire signed[31:0]    reg_activation_17_6;
wire signed[31:0]    reg_activation_17_7;
wire signed[31:0]    reg_activation_17_8;
wire signed[31:0]    reg_activation_17_9;
wire signed[31:0]    reg_activation_17_10;
wire signed[31:0]    reg_activation_17_11;
wire signed[31:0]    reg_activation_17_12;
wire signed[31:0]    reg_activation_17_13;
wire signed[31:0]    reg_activation_17_14;
wire signed[31:0]    reg_activation_17_15;
wire signed[31:0]    reg_activation_17_16;
wire signed[31:0]    reg_activation_17_17;
wire signed[31:0]    reg_activation_17_18;
wire signed[31:0]    reg_activation_17_19;
wire signed[31:0]    reg_activation_17_20;
wire signed[31:0]    reg_activation_17_21;
wire signed[31:0]    reg_activation_17_22;
wire signed[31:0]    reg_activation_17_23;
wire signed[31:0]    reg_activation_17_24;
wire signed[31:0]    reg_activation_17_25;
wire signed[31:0]    reg_activation_17_26;
wire signed[31:0]    reg_activation_17_27;
wire signed[31:0]    reg_activation_17_28;
wire signed[31:0]    reg_activation_17_29;
wire signed[31:0]    reg_activation_17_30;
wire signed[31:0]    reg_activation_17_31;
wire signed[31:0]    reg_activation_17_32;
wire signed[31:0]    reg_activation_17_33;
wire signed[31:0]    reg_activation_17_34;
wire signed[31:0]    reg_activation_17_35;
wire signed[31:0]    reg_activation_17_36;
wire signed[31:0]    reg_activation_17_37;
wire signed[31:0]    reg_activation_17_38;
wire signed[31:0]    reg_activation_17_39;
wire signed[31:0]    reg_activation_17_40;
wire signed[31:0]    reg_activation_17_41;
wire signed[31:0]    reg_activation_17_42;
wire signed[31:0]    reg_activation_17_43;
wire signed[31:0]    reg_activation_17_44;
wire signed[31:0]    reg_activation_17_45;
wire signed[31:0]    reg_activation_17_46;
wire signed[31:0]    reg_activation_17_47;
wire signed[31:0]    reg_activation_17_48;
wire signed[31:0]    reg_activation_17_49;
wire signed[31:0]    reg_activation_17_50;
wire signed[31:0]    reg_activation_17_51;
wire signed[31:0]    reg_activation_17_52;
wire signed[31:0]    reg_activation_17_53;
wire signed[31:0]    reg_activation_17_54;
wire signed[31:0]    reg_activation_17_55;
wire signed[31:0]    reg_activation_17_56;
wire signed[31:0]    reg_activation_17_57;
wire signed[31:0]    reg_activation_17_58;
wire signed[31:0]    reg_activation_17_59;
wire signed[31:0]    reg_activation_17_60;
wire signed[31:0]    reg_activation_17_61;
wire signed[31:0]    reg_activation_17_62;
wire signed[31:0]    reg_activation_17_63;
wire signed[31:0]    reg_activation_18_0;
wire signed[31:0]    reg_activation_18_1;
wire signed[31:0]    reg_activation_18_2;
wire signed[31:0]    reg_activation_18_3;
wire signed[31:0]    reg_activation_18_4;
wire signed[31:0]    reg_activation_18_5;
wire signed[31:0]    reg_activation_18_6;
wire signed[31:0]    reg_activation_18_7;
wire signed[31:0]    reg_activation_18_8;
wire signed[31:0]    reg_activation_18_9;
wire signed[31:0]    reg_activation_18_10;
wire signed[31:0]    reg_activation_18_11;
wire signed[31:0]    reg_activation_18_12;
wire signed[31:0]    reg_activation_18_13;
wire signed[31:0]    reg_activation_18_14;
wire signed[31:0]    reg_activation_18_15;
wire signed[31:0]    reg_activation_18_16;
wire signed[31:0]    reg_activation_18_17;
wire signed[31:0]    reg_activation_18_18;
wire signed[31:0]    reg_activation_18_19;
wire signed[31:0]    reg_activation_18_20;
wire signed[31:0]    reg_activation_18_21;
wire signed[31:0]    reg_activation_18_22;
wire signed[31:0]    reg_activation_18_23;
wire signed[31:0]    reg_activation_18_24;
wire signed[31:0]    reg_activation_18_25;
wire signed[31:0]    reg_activation_18_26;
wire signed[31:0]    reg_activation_18_27;
wire signed[31:0]    reg_activation_18_28;
wire signed[31:0]    reg_activation_18_29;
wire signed[31:0]    reg_activation_18_30;
wire signed[31:0]    reg_activation_18_31;
wire signed[31:0]    reg_activation_18_32;
wire signed[31:0]    reg_activation_18_33;
wire signed[31:0]    reg_activation_18_34;
wire signed[31:0]    reg_activation_18_35;
wire signed[31:0]    reg_activation_18_36;
wire signed[31:0]    reg_activation_18_37;
wire signed[31:0]    reg_activation_18_38;
wire signed[31:0]    reg_activation_18_39;
wire signed[31:0]    reg_activation_18_40;
wire signed[31:0]    reg_activation_18_41;
wire signed[31:0]    reg_activation_18_42;
wire signed[31:0]    reg_activation_18_43;
wire signed[31:0]    reg_activation_18_44;
wire signed[31:0]    reg_activation_18_45;
wire signed[31:0]    reg_activation_18_46;
wire signed[31:0]    reg_activation_18_47;
wire signed[31:0]    reg_activation_18_48;
wire signed[31:0]    reg_activation_18_49;
wire signed[31:0]    reg_activation_18_50;
wire signed[31:0]    reg_activation_18_51;
wire signed[31:0]    reg_activation_18_52;
wire signed[31:0]    reg_activation_18_53;
wire signed[31:0]    reg_activation_18_54;
wire signed[31:0]    reg_activation_18_55;
wire signed[31:0]    reg_activation_18_56;
wire signed[31:0]    reg_activation_18_57;
wire signed[31:0]    reg_activation_18_58;
wire signed[31:0]    reg_activation_18_59;
wire signed[31:0]    reg_activation_18_60;
wire signed[31:0]    reg_activation_18_61;
wire signed[31:0]    reg_activation_18_62;
wire signed[31:0]    reg_activation_18_63;
wire signed[31:0]    reg_activation_19_0;
wire signed[31:0]    reg_activation_19_1;
wire signed[31:0]    reg_activation_19_2;
wire signed[31:0]    reg_activation_19_3;
wire signed[31:0]    reg_activation_19_4;
wire signed[31:0]    reg_activation_19_5;
wire signed[31:0]    reg_activation_19_6;
wire signed[31:0]    reg_activation_19_7;
wire signed[31:0]    reg_activation_19_8;
wire signed[31:0]    reg_activation_19_9;
wire signed[31:0]    reg_activation_19_10;
wire signed[31:0]    reg_activation_19_11;
wire signed[31:0]    reg_activation_19_12;
wire signed[31:0]    reg_activation_19_13;
wire signed[31:0]    reg_activation_19_14;
wire signed[31:0]    reg_activation_19_15;
wire signed[31:0]    reg_activation_19_16;
wire signed[31:0]    reg_activation_19_17;
wire signed[31:0]    reg_activation_19_18;
wire signed[31:0]    reg_activation_19_19;
wire signed[31:0]    reg_activation_19_20;
wire signed[31:0]    reg_activation_19_21;
wire signed[31:0]    reg_activation_19_22;
wire signed[31:0]    reg_activation_19_23;
wire signed[31:0]    reg_activation_19_24;
wire signed[31:0]    reg_activation_19_25;
wire signed[31:0]    reg_activation_19_26;
wire signed[31:0]    reg_activation_19_27;
wire signed[31:0]    reg_activation_19_28;
wire signed[31:0]    reg_activation_19_29;
wire signed[31:0]    reg_activation_19_30;
wire signed[31:0]    reg_activation_19_31;
wire signed[31:0]    reg_activation_19_32;
wire signed[31:0]    reg_activation_19_33;
wire signed[31:0]    reg_activation_19_34;
wire signed[31:0]    reg_activation_19_35;
wire signed[31:0]    reg_activation_19_36;
wire signed[31:0]    reg_activation_19_37;
wire signed[31:0]    reg_activation_19_38;
wire signed[31:0]    reg_activation_19_39;
wire signed[31:0]    reg_activation_19_40;
wire signed[31:0]    reg_activation_19_41;
wire signed[31:0]    reg_activation_19_42;
wire signed[31:0]    reg_activation_19_43;
wire signed[31:0]    reg_activation_19_44;
wire signed[31:0]    reg_activation_19_45;
wire signed[31:0]    reg_activation_19_46;
wire signed[31:0]    reg_activation_19_47;
wire signed[31:0]    reg_activation_19_48;
wire signed[31:0]    reg_activation_19_49;
wire signed[31:0]    reg_activation_19_50;
wire signed[31:0]    reg_activation_19_51;
wire signed[31:0]    reg_activation_19_52;
wire signed[31:0]    reg_activation_19_53;
wire signed[31:0]    reg_activation_19_54;
wire signed[31:0]    reg_activation_19_55;
wire signed[31:0]    reg_activation_19_56;
wire signed[31:0]    reg_activation_19_57;
wire signed[31:0]    reg_activation_19_58;
wire signed[31:0]    reg_activation_19_59;
wire signed[31:0]    reg_activation_19_60;
wire signed[31:0]    reg_activation_19_61;
wire signed[31:0]    reg_activation_19_62;
wire signed[31:0]    reg_activation_19_63;
wire signed[31:0]    reg_activation_20_0;
wire signed[31:0]    reg_activation_20_1;
wire signed[31:0]    reg_activation_20_2;
wire signed[31:0]    reg_activation_20_3;
wire signed[31:0]    reg_activation_20_4;
wire signed[31:0]    reg_activation_20_5;
wire signed[31:0]    reg_activation_20_6;
wire signed[31:0]    reg_activation_20_7;
wire signed[31:0]    reg_activation_20_8;
wire signed[31:0]    reg_activation_20_9;
wire signed[31:0]    reg_activation_20_10;
wire signed[31:0]    reg_activation_20_11;
wire signed[31:0]    reg_activation_20_12;
wire signed[31:0]    reg_activation_20_13;
wire signed[31:0]    reg_activation_20_14;
wire signed[31:0]    reg_activation_20_15;
wire signed[31:0]    reg_activation_20_16;
wire signed[31:0]    reg_activation_20_17;
wire signed[31:0]    reg_activation_20_18;
wire signed[31:0]    reg_activation_20_19;
wire signed[31:0]    reg_activation_20_20;
wire signed[31:0]    reg_activation_20_21;
wire signed[31:0]    reg_activation_20_22;
wire signed[31:0]    reg_activation_20_23;
wire signed[31:0]    reg_activation_20_24;
wire signed[31:0]    reg_activation_20_25;
wire signed[31:0]    reg_activation_20_26;
wire signed[31:0]    reg_activation_20_27;
wire signed[31:0]    reg_activation_20_28;
wire signed[31:0]    reg_activation_20_29;
wire signed[31:0]    reg_activation_20_30;
wire signed[31:0]    reg_activation_20_31;
wire signed[31:0]    reg_activation_20_32;
wire signed[31:0]    reg_activation_20_33;
wire signed[31:0]    reg_activation_20_34;
wire signed[31:0]    reg_activation_20_35;
wire signed[31:0]    reg_activation_20_36;
wire signed[31:0]    reg_activation_20_37;
wire signed[31:0]    reg_activation_20_38;
wire signed[31:0]    reg_activation_20_39;
wire signed[31:0]    reg_activation_20_40;
wire signed[31:0]    reg_activation_20_41;
wire signed[31:0]    reg_activation_20_42;
wire signed[31:0]    reg_activation_20_43;
wire signed[31:0]    reg_activation_20_44;
wire signed[31:0]    reg_activation_20_45;
wire signed[31:0]    reg_activation_20_46;
wire signed[31:0]    reg_activation_20_47;
wire signed[31:0]    reg_activation_20_48;
wire signed[31:0]    reg_activation_20_49;
wire signed[31:0]    reg_activation_20_50;
wire signed[31:0]    reg_activation_20_51;
wire signed[31:0]    reg_activation_20_52;
wire signed[31:0]    reg_activation_20_53;
wire signed[31:0]    reg_activation_20_54;
wire signed[31:0]    reg_activation_20_55;
wire signed[31:0]    reg_activation_20_56;
wire signed[31:0]    reg_activation_20_57;
wire signed[31:0]    reg_activation_20_58;
wire signed[31:0]    reg_activation_20_59;
wire signed[31:0]    reg_activation_20_60;
wire signed[31:0]    reg_activation_20_61;
wire signed[31:0]    reg_activation_20_62;
wire signed[31:0]    reg_activation_20_63;
wire signed[31:0]    reg_activation_21_0;
wire signed[31:0]    reg_activation_21_1;
wire signed[31:0]    reg_activation_21_2;
wire signed[31:0]    reg_activation_21_3;
wire signed[31:0]    reg_activation_21_4;
wire signed[31:0]    reg_activation_21_5;
wire signed[31:0]    reg_activation_21_6;
wire signed[31:0]    reg_activation_21_7;
wire signed[31:0]    reg_activation_21_8;
wire signed[31:0]    reg_activation_21_9;
wire signed[31:0]    reg_activation_21_10;
wire signed[31:0]    reg_activation_21_11;
wire signed[31:0]    reg_activation_21_12;
wire signed[31:0]    reg_activation_21_13;
wire signed[31:0]    reg_activation_21_14;
wire signed[31:0]    reg_activation_21_15;
wire signed[31:0]    reg_activation_21_16;
wire signed[31:0]    reg_activation_21_17;
wire signed[31:0]    reg_activation_21_18;
wire signed[31:0]    reg_activation_21_19;
wire signed[31:0]    reg_activation_21_20;
wire signed[31:0]    reg_activation_21_21;
wire signed[31:0]    reg_activation_21_22;
wire signed[31:0]    reg_activation_21_23;
wire signed[31:0]    reg_activation_21_24;
wire signed[31:0]    reg_activation_21_25;
wire signed[31:0]    reg_activation_21_26;
wire signed[31:0]    reg_activation_21_27;
wire signed[31:0]    reg_activation_21_28;
wire signed[31:0]    reg_activation_21_29;
wire signed[31:0]    reg_activation_21_30;
wire signed[31:0]    reg_activation_21_31;
wire signed[31:0]    reg_activation_21_32;
wire signed[31:0]    reg_activation_21_33;
wire signed[31:0]    reg_activation_21_34;
wire signed[31:0]    reg_activation_21_35;
wire signed[31:0]    reg_activation_21_36;
wire signed[31:0]    reg_activation_21_37;
wire signed[31:0]    reg_activation_21_38;
wire signed[31:0]    reg_activation_21_39;
wire signed[31:0]    reg_activation_21_40;
wire signed[31:0]    reg_activation_21_41;
wire signed[31:0]    reg_activation_21_42;
wire signed[31:0]    reg_activation_21_43;
wire signed[31:0]    reg_activation_21_44;
wire signed[31:0]    reg_activation_21_45;
wire signed[31:0]    reg_activation_21_46;
wire signed[31:0]    reg_activation_21_47;
wire signed[31:0]    reg_activation_21_48;
wire signed[31:0]    reg_activation_21_49;
wire signed[31:0]    reg_activation_21_50;
wire signed[31:0]    reg_activation_21_51;
wire signed[31:0]    reg_activation_21_52;
wire signed[31:0]    reg_activation_21_53;
wire signed[31:0]    reg_activation_21_54;
wire signed[31:0]    reg_activation_21_55;
wire signed[31:0]    reg_activation_21_56;
wire signed[31:0]    reg_activation_21_57;
wire signed[31:0]    reg_activation_21_58;
wire signed[31:0]    reg_activation_21_59;
wire signed[31:0]    reg_activation_21_60;
wire signed[31:0]    reg_activation_21_61;
wire signed[31:0]    reg_activation_21_62;
wire signed[31:0]    reg_activation_21_63;
wire signed[31:0]    reg_activation_22_0;
wire signed[31:0]    reg_activation_22_1;
wire signed[31:0]    reg_activation_22_2;
wire signed[31:0]    reg_activation_22_3;
wire signed[31:0]    reg_activation_22_4;
wire signed[31:0]    reg_activation_22_5;
wire signed[31:0]    reg_activation_22_6;
wire signed[31:0]    reg_activation_22_7;
wire signed[31:0]    reg_activation_22_8;
wire signed[31:0]    reg_activation_22_9;
wire signed[31:0]    reg_activation_22_10;
wire signed[31:0]    reg_activation_22_11;
wire signed[31:0]    reg_activation_22_12;
wire signed[31:0]    reg_activation_22_13;
wire signed[31:0]    reg_activation_22_14;
wire signed[31:0]    reg_activation_22_15;
wire signed[31:0]    reg_activation_22_16;
wire signed[31:0]    reg_activation_22_17;
wire signed[31:0]    reg_activation_22_18;
wire signed[31:0]    reg_activation_22_19;
wire signed[31:0]    reg_activation_22_20;
wire signed[31:0]    reg_activation_22_21;
wire signed[31:0]    reg_activation_22_22;
wire signed[31:0]    reg_activation_22_23;
wire signed[31:0]    reg_activation_22_24;
wire signed[31:0]    reg_activation_22_25;
wire signed[31:0]    reg_activation_22_26;
wire signed[31:0]    reg_activation_22_27;
wire signed[31:0]    reg_activation_22_28;
wire signed[31:0]    reg_activation_22_29;
wire signed[31:0]    reg_activation_22_30;
wire signed[31:0]    reg_activation_22_31;
wire signed[31:0]    reg_activation_22_32;
wire signed[31:0]    reg_activation_22_33;
wire signed[31:0]    reg_activation_22_34;
wire signed[31:0]    reg_activation_22_35;
wire signed[31:0]    reg_activation_22_36;
wire signed[31:0]    reg_activation_22_37;
wire signed[31:0]    reg_activation_22_38;
wire signed[31:0]    reg_activation_22_39;
wire signed[31:0]    reg_activation_22_40;
wire signed[31:0]    reg_activation_22_41;
wire signed[31:0]    reg_activation_22_42;
wire signed[31:0]    reg_activation_22_43;
wire signed[31:0]    reg_activation_22_44;
wire signed[31:0]    reg_activation_22_45;
wire signed[31:0]    reg_activation_22_46;
wire signed[31:0]    reg_activation_22_47;
wire signed[31:0]    reg_activation_22_48;
wire signed[31:0]    reg_activation_22_49;
wire signed[31:0]    reg_activation_22_50;
wire signed[31:0]    reg_activation_22_51;
wire signed[31:0]    reg_activation_22_52;
wire signed[31:0]    reg_activation_22_53;
wire signed[31:0]    reg_activation_22_54;
wire signed[31:0]    reg_activation_22_55;
wire signed[31:0]    reg_activation_22_56;
wire signed[31:0]    reg_activation_22_57;
wire signed[31:0]    reg_activation_22_58;
wire signed[31:0]    reg_activation_22_59;
wire signed[31:0]    reg_activation_22_60;
wire signed[31:0]    reg_activation_22_61;
wire signed[31:0]    reg_activation_22_62;
wire signed[31:0]    reg_activation_22_63;
wire signed[31:0]    reg_activation_23_0;
wire signed[31:0]    reg_activation_23_1;
wire signed[31:0]    reg_activation_23_2;
wire signed[31:0]    reg_activation_23_3;
wire signed[31:0]    reg_activation_23_4;
wire signed[31:0]    reg_activation_23_5;
wire signed[31:0]    reg_activation_23_6;
wire signed[31:0]    reg_activation_23_7;
wire signed[31:0]    reg_activation_23_8;
wire signed[31:0]    reg_activation_23_9;
wire signed[31:0]    reg_activation_23_10;
wire signed[31:0]    reg_activation_23_11;
wire signed[31:0]    reg_activation_23_12;
wire signed[31:0]    reg_activation_23_13;
wire signed[31:0]    reg_activation_23_14;
wire signed[31:0]    reg_activation_23_15;
wire signed[31:0]    reg_activation_23_16;
wire signed[31:0]    reg_activation_23_17;
wire signed[31:0]    reg_activation_23_18;
wire signed[31:0]    reg_activation_23_19;
wire signed[31:0]    reg_activation_23_20;
wire signed[31:0]    reg_activation_23_21;
wire signed[31:0]    reg_activation_23_22;
wire signed[31:0]    reg_activation_23_23;
wire signed[31:0]    reg_activation_23_24;
wire signed[31:0]    reg_activation_23_25;
wire signed[31:0]    reg_activation_23_26;
wire signed[31:0]    reg_activation_23_27;
wire signed[31:0]    reg_activation_23_28;
wire signed[31:0]    reg_activation_23_29;
wire signed[31:0]    reg_activation_23_30;
wire signed[31:0]    reg_activation_23_31;
wire signed[31:0]    reg_activation_23_32;
wire signed[31:0]    reg_activation_23_33;
wire signed[31:0]    reg_activation_23_34;
wire signed[31:0]    reg_activation_23_35;
wire signed[31:0]    reg_activation_23_36;
wire signed[31:0]    reg_activation_23_37;
wire signed[31:0]    reg_activation_23_38;
wire signed[31:0]    reg_activation_23_39;
wire signed[31:0]    reg_activation_23_40;
wire signed[31:0]    reg_activation_23_41;
wire signed[31:0]    reg_activation_23_42;
wire signed[31:0]    reg_activation_23_43;
wire signed[31:0]    reg_activation_23_44;
wire signed[31:0]    reg_activation_23_45;
wire signed[31:0]    reg_activation_23_46;
wire signed[31:0]    reg_activation_23_47;
wire signed[31:0]    reg_activation_23_48;
wire signed[31:0]    reg_activation_23_49;
wire signed[31:0]    reg_activation_23_50;
wire signed[31:0]    reg_activation_23_51;
wire signed[31:0]    reg_activation_23_52;
wire signed[31:0]    reg_activation_23_53;
wire signed[31:0]    reg_activation_23_54;
wire signed[31:0]    reg_activation_23_55;
wire signed[31:0]    reg_activation_23_56;
wire signed[31:0]    reg_activation_23_57;
wire signed[31:0]    reg_activation_23_58;
wire signed[31:0]    reg_activation_23_59;
wire signed[31:0]    reg_activation_23_60;
wire signed[31:0]    reg_activation_23_61;
wire signed[31:0]    reg_activation_23_62;
wire signed[31:0]    reg_activation_23_63;
wire signed[31:0]    reg_activation_24_0;
wire signed[31:0]    reg_activation_24_1;
wire signed[31:0]    reg_activation_24_2;
wire signed[31:0]    reg_activation_24_3;
wire signed[31:0]    reg_activation_24_4;
wire signed[31:0]    reg_activation_24_5;
wire signed[31:0]    reg_activation_24_6;
wire signed[31:0]    reg_activation_24_7;
wire signed[31:0]    reg_activation_24_8;
wire signed[31:0]    reg_activation_24_9;
wire signed[31:0]    reg_activation_24_10;
wire signed[31:0]    reg_activation_24_11;
wire signed[31:0]    reg_activation_24_12;
wire signed[31:0]    reg_activation_24_13;
wire signed[31:0]    reg_activation_24_14;
wire signed[31:0]    reg_activation_24_15;
wire signed[31:0]    reg_activation_24_16;
wire signed[31:0]    reg_activation_24_17;
wire signed[31:0]    reg_activation_24_18;
wire signed[31:0]    reg_activation_24_19;
wire signed[31:0]    reg_activation_24_20;
wire signed[31:0]    reg_activation_24_21;
wire signed[31:0]    reg_activation_24_22;
wire signed[31:0]    reg_activation_24_23;
wire signed[31:0]    reg_activation_24_24;
wire signed[31:0]    reg_activation_24_25;
wire signed[31:0]    reg_activation_24_26;
wire signed[31:0]    reg_activation_24_27;
wire signed[31:0]    reg_activation_24_28;
wire signed[31:0]    reg_activation_24_29;
wire signed[31:0]    reg_activation_24_30;
wire signed[31:0]    reg_activation_24_31;
wire signed[31:0]    reg_activation_24_32;
wire signed[31:0]    reg_activation_24_33;
wire signed[31:0]    reg_activation_24_34;
wire signed[31:0]    reg_activation_24_35;
wire signed[31:0]    reg_activation_24_36;
wire signed[31:0]    reg_activation_24_37;
wire signed[31:0]    reg_activation_24_38;
wire signed[31:0]    reg_activation_24_39;
wire signed[31:0]    reg_activation_24_40;
wire signed[31:0]    reg_activation_24_41;
wire signed[31:0]    reg_activation_24_42;
wire signed[31:0]    reg_activation_24_43;
wire signed[31:0]    reg_activation_24_44;
wire signed[31:0]    reg_activation_24_45;
wire signed[31:0]    reg_activation_24_46;
wire signed[31:0]    reg_activation_24_47;
wire signed[31:0]    reg_activation_24_48;
wire signed[31:0]    reg_activation_24_49;
wire signed[31:0]    reg_activation_24_50;
wire signed[31:0]    reg_activation_24_51;
wire signed[31:0]    reg_activation_24_52;
wire signed[31:0]    reg_activation_24_53;
wire signed[31:0]    reg_activation_24_54;
wire signed[31:0]    reg_activation_24_55;
wire signed[31:0]    reg_activation_24_56;
wire signed[31:0]    reg_activation_24_57;
wire signed[31:0]    reg_activation_24_58;
wire signed[31:0]    reg_activation_24_59;
wire signed[31:0]    reg_activation_24_60;
wire signed[31:0]    reg_activation_24_61;
wire signed[31:0]    reg_activation_24_62;
wire signed[31:0]    reg_activation_24_63;
wire signed[31:0]    reg_activation_25_0;
wire signed[31:0]    reg_activation_25_1;
wire signed[31:0]    reg_activation_25_2;
wire signed[31:0]    reg_activation_25_3;
wire signed[31:0]    reg_activation_25_4;
wire signed[31:0]    reg_activation_25_5;
wire signed[31:0]    reg_activation_25_6;
wire signed[31:0]    reg_activation_25_7;
wire signed[31:0]    reg_activation_25_8;
wire signed[31:0]    reg_activation_25_9;
wire signed[31:0]    reg_activation_25_10;
wire signed[31:0]    reg_activation_25_11;
wire signed[31:0]    reg_activation_25_12;
wire signed[31:0]    reg_activation_25_13;
wire signed[31:0]    reg_activation_25_14;
wire signed[31:0]    reg_activation_25_15;
wire signed[31:0]    reg_activation_25_16;
wire signed[31:0]    reg_activation_25_17;
wire signed[31:0]    reg_activation_25_18;
wire signed[31:0]    reg_activation_25_19;
wire signed[31:0]    reg_activation_25_20;
wire signed[31:0]    reg_activation_25_21;
wire signed[31:0]    reg_activation_25_22;
wire signed[31:0]    reg_activation_25_23;
wire signed[31:0]    reg_activation_25_24;
wire signed[31:0]    reg_activation_25_25;
wire signed[31:0]    reg_activation_25_26;
wire signed[31:0]    reg_activation_25_27;
wire signed[31:0]    reg_activation_25_28;
wire signed[31:0]    reg_activation_25_29;
wire signed[31:0]    reg_activation_25_30;
wire signed[31:0]    reg_activation_25_31;
wire signed[31:0]    reg_activation_25_32;
wire signed[31:0]    reg_activation_25_33;
wire signed[31:0]    reg_activation_25_34;
wire signed[31:0]    reg_activation_25_35;
wire signed[31:0]    reg_activation_25_36;
wire signed[31:0]    reg_activation_25_37;
wire signed[31:0]    reg_activation_25_38;
wire signed[31:0]    reg_activation_25_39;
wire signed[31:0]    reg_activation_25_40;
wire signed[31:0]    reg_activation_25_41;
wire signed[31:0]    reg_activation_25_42;
wire signed[31:0]    reg_activation_25_43;
wire signed[31:0]    reg_activation_25_44;
wire signed[31:0]    reg_activation_25_45;
wire signed[31:0]    reg_activation_25_46;
wire signed[31:0]    reg_activation_25_47;
wire signed[31:0]    reg_activation_25_48;
wire signed[31:0]    reg_activation_25_49;
wire signed[31:0]    reg_activation_25_50;
wire signed[31:0]    reg_activation_25_51;
wire signed[31:0]    reg_activation_25_52;
wire signed[31:0]    reg_activation_25_53;
wire signed[31:0]    reg_activation_25_54;
wire signed[31:0]    reg_activation_25_55;
wire signed[31:0]    reg_activation_25_56;
wire signed[31:0]    reg_activation_25_57;
wire signed[31:0]    reg_activation_25_58;
wire signed[31:0]    reg_activation_25_59;
wire signed[31:0]    reg_activation_25_60;
wire signed[31:0]    reg_activation_25_61;
wire signed[31:0]    reg_activation_25_62;
wire signed[31:0]    reg_activation_25_63;
wire signed[31:0]    reg_activation_26_0;
wire signed[31:0]    reg_activation_26_1;
wire signed[31:0]    reg_activation_26_2;
wire signed[31:0]    reg_activation_26_3;
wire signed[31:0]    reg_activation_26_4;
wire signed[31:0]    reg_activation_26_5;
wire signed[31:0]    reg_activation_26_6;
wire signed[31:0]    reg_activation_26_7;
wire signed[31:0]    reg_activation_26_8;
wire signed[31:0]    reg_activation_26_9;
wire signed[31:0]    reg_activation_26_10;
wire signed[31:0]    reg_activation_26_11;
wire signed[31:0]    reg_activation_26_12;
wire signed[31:0]    reg_activation_26_13;
wire signed[31:0]    reg_activation_26_14;
wire signed[31:0]    reg_activation_26_15;
wire signed[31:0]    reg_activation_26_16;
wire signed[31:0]    reg_activation_26_17;
wire signed[31:0]    reg_activation_26_18;
wire signed[31:0]    reg_activation_26_19;
wire signed[31:0]    reg_activation_26_20;
wire signed[31:0]    reg_activation_26_21;
wire signed[31:0]    reg_activation_26_22;
wire signed[31:0]    reg_activation_26_23;
wire signed[31:0]    reg_activation_26_24;
wire signed[31:0]    reg_activation_26_25;
wire signed[31:0]    reg_activation_26_26;
wire signed[31:0]    reg_activation_26_27;
wire signed[31:0]    reg_activation_26_28;
wire signed[31:0]    reg_activation_26_29;
wire signed[31:0]    reg_activation_26_30;
wire signed[31:0]    reg_activation_26_31;
wire signed[31:0]    reg_activation_26_32;
wire signed[31:0]    reg_activation_26_33;
wire signed[31:0]    reg_activation_26_34;
wire signed[31:0]    reg_activation_26_35;
wire signed[31:0]    reg_activation_26_36;
wire signed[31:0]    reg_activation_26_37;
wire signed[31:0]    reg_activation_26_38;
wire signed[31:0]    reg_activation_26_39;
wire signed[31:0]    reg_activation_26_40;
wire signed[31:0]    reg_activation_26_41;
wire signed[31:0]    reg_activation_26_42;
wire signed[31:0]    reg_activation_26_43;
wire signed[31:0]    reg_activation_26_44;
wire signed[31:0]    reg_activation_26_45;
wire signed[31:0]    reg_activation_26_46;
wire signed[31:0]    reg_activation_26_47;
wire signed[31:0]    reg_activation_26_48;
wire signed[31:0]    reg_activation_26_49;
wire signed[31:0]    reg_activation_26_50;
wire signed[31:0]    reg_activation_26_51;
wire signed[31:0]    reg_activation_26_52;
wire signed[31:0]    reg_activation_26_53;
wire signed[31:0]    reg_activation_26_54;
wire signed[31:0]    reg_activation_26_55;
wire signed[31:0]    reg_activation_26_56;
wire signed[31:0]    reg_activation_26_57;
wire signed[31:0]    reg_activation_26_58;
wire signed[31:0]    reg_activation_26_59;
wire signed[31:0]    reg_activation_26_60;
wire signed[31:0]    reg_activation_26_61;
wire signed[31:0]    reg_activation_26_62;
wire signed[31:0]    reg_activation_26_63;
wire signed[31:0]    reg_activation_27_0;
wire signed[31:0]    reg_activation_27_1;
wire signed[31:0]    reg_activation_27_2;
wire signed[31:0]    reg_activation_27_3;
wire signed[31:0]    reg_activation_27_4;
wire signed[31:0]    reg_activation_27_5;
wire signed[31:0]    reg_activation_27_6;
wire signed[31:0]    reg_activation_27_7;
wire signed[31:0]    reg_activation_27_8;
wire signed[31:0]    reg_activation_27_9;
wire signed[31:0]    reg_activation_27_10;
wire signed[31:0]    reg_activation_27_11;
wire signed[31:0]    reg_activation_27_12;
wire signed[31:0]    reg_activation_27_13;
wire signed[31:0]    reg_activation_27_14;
wire signed[31:0]    reg_activation_27_15;
wire signed[31:0]    reg_activation_27_16;
wire signed[31:0]    reg_activation_27_17;
wire signed[31:0]    reg_activation_27_18;
wire signed[31:0]    reg_activation_27_19;
wire signed[31:0]    reg_activation_27_20;
wire signed[31:0]    reg_activation_27_21;
wire signed[31:0]    reg_activation_27_22;
wire signed[31:0]    reg_activation_27_23;
wire signed[31:0]    reg_activation_27_24;
wire signed[31:0]    reg_activation_27_25;
wire signed[31:0]    reg_activation_27_26;
wire signed[31:0]    reg_activation_27_27;
wire signed[31:0]    reg_activation_27_28;
wire signed[31:0]    reg_activation_27_29;
wire signed[31:0]    reg_activation_27_30;
wire signed[31:0]    reg_activation_27_31;
wire signed[31:0]    reg_activation_27_32;
wire signed[31:0]    reg_activation_27_33;
wire signed[31:0]    reg_activation_27_34;
wire signed[31:0]    reg_activation_27_35;
wire signed[31:0]    reg_activation_27_36;
wire signed[31:0]    reg_activation_27_37;
wire signed[31:0]    reg_activation_27_38;
wire signed[31:0]    reg_activation_27_39;
wire signed[31:0]    reg_activation_27_40;
wire signed[31:0]    reg_activation_27_41;
wire signed[31:0]    reg_activation_27_42;
wire signed[31:0]    reg_activation_27_43;
wire signed[31:0]    reg_activation_27_44;
wire signed[31:0]    reg_activation_27_45;
wire signed[31:0]    reg_activation_27_46;
wire signed[31:0]    reg_activation_27_47;
wire signed[31:0]    reg_activation_27_48;
wire signed[31:0]    reg_activation_27_49;
wire signed[31:0]    reg_activation_27_50;
wire signed[31:0]    reg_activation_27_51;
wire signed[31:0]    reg_activation_27_52;
wire signed[31:0]    reg_activation_27_53;
wire signed[31:0]    reg_activation_27_54;
wire signed[31:0]    reg_activation_27_55;
wire signed[31:0]    reg_activation_27_56;
wire signed[31:0]    reg_activation_27_57;
wire signed[31:0]    reg_activation_27_58;
wire signed[31:0]    reg_activation_27_59;
wire signed[31:0]    reg_activation_27_60;
wire signed[31:0]    reg_activation_27_61;
wire signed[31:0]    reg_activation_27_62;
wire signed[31:0]    reg_activation_27_63;
wire signed[31:0]    reg_activation_28_0;
wire signed[31:0]    reg_activation_28_1;
wire signed[31:0]    reg_activation_28_2;
wire signed[31:0]    reg_activation_28_3;
wire signed[31:0]    reg_activation_28_4;
wire signed[31:0]    reg_activation_28_5;
wire signed[31:0]    reg_activation_28_6;
wire signed[31:0]    reg_activation_28_7;
wire signed[31:0]    reg_activation_28_8;
wire signed[31:0]    reg_activation_28_9;
wire signed[31:0]    reg_activation_28_10;
wire signed[31:0]    reg_activation_28_11;
wire signed[31:0]    reg_activation_28_12;
wire signed[31:0]    reg_activation_28_13;
wire signed[31:0]    reg_activation_28_14;
wire signed[31:0]    reg_activation_28_15;
wire signed[31:0]    reg_activation_28_16;
wire signed[31:0]    reg_activation_28_17;
wire signed[31:0]    reg_activation_28_18;
wire signed[31:0]    reg_activation_28_19;
wire signed[31:0]    reg_activation_28_20;
wire signed[31:0]    reg_activation_28_21;
wire signed[31:0]    reg_activation_28_22;
wire signed[31:0]    reg_activation_28_23;
wire signed[31:0]    reg_activation_28_24;
wire signed[31:0]    reg_activation_28_25;
wire signed[31:0]    reg_activation_28_26;
wire signed[31:0]    reg_activation_28_27;
wire signed[31:0]    reg_activation_28_28;
wire signed[31:0]    reg_activation_28_29;
wire signed[31:0]    reg_activation_28_30;
wire signed[31:0]    reg_activation_28_31;
wire signed[31:0]    reg_activation_28_32;
wire signed[31:0]    reg_activation_28_33;
wire signed[31:0]    reg_activation_28_34;
wire signed[31:0]    reg_activation_28_35;
wire signed[31:0]    reg_activation_28_36;
wire signed[31:0]    reg_activation_28_37;
wire signed[31:0]    reg_activation_28_38;
wire signed[31:0]    reg_activation_28_39;
wire signed[31:0]    reg_activation_28_40;
wire signed[31:0]    reg_activation_28_41;
wire signed[31:0]    reg_activation_28_42;
wire signed[31:0]    reg_activation_28_43;
wire signed[31:0]    reg_activation_28_44;
wire signed[31:0]    reg_activation_28_45;
wire signed[31:0]    reg_activation_28_46;
wire signed[31:0]    reg_activation_28_47;
wire signed[31:0]    reg_activation_28_48;
wire signed[31:0]    reg_activation_28_49;
wire signed[31:0]    reg_activation_28_50;
wire signed[31:0]    reg_activation_28_51;
wire signed[31:0]    reg_activation_28_52;
wire signed[31:0]    reg_activation_28_53;
wire signed[31:0]    reg_activation_28_54;
wire signed[31:0]    reg_activation_28_55;
wire signed[31:0]    reg_activation_28_56;
wire signed[31:0]    reg_activation_28_57;
wire signed[31:0]    reg_activation_28_58;
wire signed[31:0]    reg_activation_28_59;
wire signed[31:0]    reg_activation_28_60;
wire signed[31:0]    reg_activation_28_61;
wire signed[31:0]    reg_activation_28_62;
wire signed[31:0]    reg_activation_28_63;
wire signed[31:0]    reg_activation_29_0;
wire signed[31:0]    reg_activation_29_1;
wire signed[31:0]    reg_activation_29_2;
wire signed[31:0]    reg_activation_29_3;
wire signed[31:0]    reg_activation_29_4;
wire signed[31:0]    reg_activation_29_5;
wire signed[31:0]    reg_activation_29_6;
wire signed[31:0]    reg_activation_29_7;
wire signed[31:0]    reg_activation_29_8;
wire signed[31:0]    reg_activation_29_9;
wire signed[31:0]    reg_activation_29_10;
wire signed[31:0]    reg_activation_29_11;
wire signed[31:0]    reg_activation_29_12;
wire signed[31:0]    reg_activation_29_13;
wire signed[31:0]    reg_activation_29_14;
wire signed[31:0]    reg_activation_29_15;
wire signed[31:0]    reg_activation_29_16;
wire signed[31:0]    reg_activation_29_17;
wire signed[31:0]    reg_activation_29_18;
wire signed[31:0]    reg_activation_29_19;
wire signed[31:0]    reg_activation_29_20;
wire signed[31:0]    reg_activation_29_21;
wire signed[31:0]    reg_activation_29_22;
wire signed[31:0]    reg_activation_29_23;
wire signed[31:0]    reg_activation_29_24;
wire signed[31:0]    reg_activation_29_25;
wire signed[31:0]    reg_activation_29_26;
wire signed[31:0]    reg_activation_29_27;
wire signed[31:0]    reg_activation_29_28;
wire signed[31:0]    reg_activation_29_29;
wire signed[31:0]    reg_activation_29_30;
wire signed[31:0]    reg_activation_29_31;
wire signed[31:0]    reg_activation_29_32;
wire signed[31:0]    reg_activation_29_33;
wire signed[31:0]    reg_activation_29_34;
wire signed[31:0]    reg_activation_29_35;
wire signed[31:0]    reg_activation_29_36;
wire signed[31:0]    reg_activation_29_37;
wire signed[31:0]    reg_activation_29_38;
wire signed[31:0]    reg_activation_29_39;
wire signed[31:0]    reg_activation_29_40;
wire signed[31:0]    reg_activation_29_41;
wire signed[31:0]    reg_activation_29_42;
wire signed[31:0]    reg_activation_29_43;
wire signed[31:0]    reg_activation_29_44;
wire signed[31:0]    reg_activation_29_45;
wire signed[31:0]    reg_activation_29_46;
wire signed[31:0]    reg_activation_29_47;
wire signed[31:0]    reg_activation_29_48;
wire signed[31:0]    reg_activation_29_49;
wire signed[31:0]    reg_activation_29_50;
wire signed[31:0]    reg_activation_29_51;
wire signed[31:0]    reg_activation_29_52;
wire signed[31:0]    reg_activation_29_53;
wire signed[31:0]    reg_activation_29_54;
wire signed[31:0]    reg_activation_29_55;
wire signed[31:0]    reg_activation_29_56;
wire signed[31:0]    reg_activation_29_57;
wire signed[31:0]    reg_activation_29_58;
wire signed[31:0]    reg_activation_29_59;
wire signed[31:0]    reg_activation_29_60;
wire signed[31:0]    reg_activation_29_61;
wire signed[31:0]    reg_activation_29_62;
wire signed[31:0]    reg_activation_29_63;
wire signed[31:0]    reg_activation_30_0;
wire signed[31:0]    reg_activation_30_1;
wire signed[31:0]    reg_activation_30_2;
wire signed[31:0]    reg_activation_30_3;
wire signed[31:0]    reg_activation_30_4;
wire signed[31:0]    reg_activation_30_5;
wire signed[31:0]    reg_activation_30_6;
wire signed[31:0]    reg_activation_30_7;
wire signed[31:0]    reg_activation_30_8;
wire signed[31:0]    reg_activation_30_9;
wire signed[31:0]    reg_activation_30_10;
wire signed[31:0]    reg_activation_30_11;
wire signed[31:0]    reg_activation_30_12;
wire signed[31:0]    reg_activation_30_13;
wire signed[31:0]    reg_activation_30_14;
wire signed[31:0]    reg_activation_30_15;
wire signed[31:0]    reg_activation_30_16;
wire signed[31:0]    reg_activation_30_17;
wire signed[31:0]    reg_activation_30_18;
wire signed[31:0]    reg_activation_30_19;
wire signed[31:0]    reg_activation_30_20;
wire signed[31:0]    reg_activation_30_21;
wire signed[31:0]    reg_activation_30_22;
wire signed[31:0]    reg_activation_30_23;
wire signed[31:0]    reg_activation_30_24;
wire signed[31:0]    reg_activation_30_25;
wire signed[31:0]    reg_activation_30_26;
wire signed[31:0]    reg_activation_30_27;
wire signed[31:0]    reg_activation_30_28;
wire signed[31:0]    reg_activation_30_29;
wire signed[31:0]    reg_activation_30_30;
wire signed[31:0]    reg_activation_30_31;
wire signed[31:0]    reg_activation_30_32;
wire signed[31:0]    reg_activation_30_33;
wire signed[31:0]    reg_activation_30_34;
wire signed[31:0]    reg_activation_30_35;
wire signed[31:0]    reg_activation_30_36;
wire signed[31:0]    reg_activation_30_37;
wire signed[31:0]    reg_activation_30_38;
wire signed[31:0]    reg_activation_30_39;
wire signed[31:0]    reg_activation_30_40;
wire signed[31:0]    reg_activation_30_41;
wire signed[31:0]    reg_activation_30_42;
wire signed[31:0]    reg_activation_30_43;
wire signed[31:0]    reg_activation_30_44;
wire signed[31:0]    reg_activation_30_45;
wire signed[31:0]    reg_activation_30_46;
wire signed[31:0]    reg_activation_30_47;
wire signed[31:0]    reg_activation_30_48;
wire signed[31:0]    reg_activation_30_49;
wire signed[31:0]    reg_activation_30_50;
wire signed[31:0]    reg_activation_30_51;
wire signed[31:0]    reg_activation_30_52;
wire signed[31:0]    reg_activation_30_53;
wire signed[31:0]    reg_activation_30_54;
wire signed[31:0]    reg_activation_30_55;
wire signed[31:0]    reg_activation_30_56;
wire signed[31:0]    reg_activation_30_57;
wire signed[31:0]    reg_activation_30_58;
wire signed[31:0]    reg_activation_30_59;
wire signed[31:0]    reg_activation_30_60;
wire signed[31:0]    reg_activation_30_61;
wire signed[31:0]    reg_activation_30_62;
wire signed[31:0]    reg_activation_30_63;
wire signed[31:0]    reg_activation_31_0;
wire signed[31:0]    reg_activation_31_1;
wire signed[31:0]    reg_activation_31_2;
wire signed[31:0]    reg_activation_31_3;
wire signed[31:0]    reg_activation_31_4;
wire signed[31:0]    reg_activation_31_5;
wire signed[31:0]    reg_activation_31_6;
wire signed[31:0]    reg_activation_31_7;
wire signed[31:0]    reg_activation_31_8;
wire signed[31:0]    reg_activation_31_9;
wire signed[31:0]    reg_activation_31_10;
wire signed[31:0]    reg_activation_31_11;
wire signed[31:0]    reg_activation_31_12;
wire signed[31:0]    reg_activation_31_13;
wire signed[31:0]    reg_activation_31_14;
wire signed[31:0]    reg_activation_31_15;
wire signed[31:0]    reg_activation_31_16;
wire signed[31:0]    reg_activation_31_17;
wire signed[31:0]    reg_activation_31_18;
wire signed[31:0]    reg_activation_31_19;
wire signed[31:0]    reg_activation_31_20;
wire signed[31:0]    reg_activation_31_21;
wire signed[31:0]    reg_activation_31_22;
wire signed[31:0]    reg_activation_31_23;
wire signed[31:0]    reg_activation_31_24;
wire signed[31:0]    reg_activation_31_25;
wire signed[31:0]    reg_activation_31_26;
wire signed[31:0]    reg_activation_31_27;
wire signed[31:0]    reg_activation_31_28;
wire signed[31:0]    reg_activation_31_29;
wire signed[31:0]    reg_activation_31_30;
wire signed[31:0]    reg_activation_31_31;
wire signed[31:0]    reg_activation_31_32;
wire signed[31:0]    reg_activation_31_33;
wire signed[31:0]    reg_activation_31_34;
wire signed[31:0]    reg_activation_31_35;
wire signed[31:0]    reg_activation_31_36;
wire signed[31:0]    reg_activation_31_37;
wire signed[31:0]    reg_activation_31_38;
wire signed[31:0]    reg_activation_31_39;
wire signed[31:0]    reg_activation_31_40;
wire signed[31:0]    reg_activation_31_41;
wire signed[31:0]    reg_activation_31_42;
wire signed[31:0]    reg_activation_31_43;
wire signed[31:0]    reg_activation_31_44;
wire signed[31:0]    reg_activation_31_45;
wire signed[31:0]    reg_activation_31_46;
wire signed[31:0]    reg_activation_31_47;
wire signed[31:0]    reg_activation_31_48;
wire signed[31:0]    reg_activation_31_49;
wire signed[31:0]    reg_activation_31_50;
wire signed[31:0]    reg_activation_31_51;
wire signed[31:0]    reg_activation_31_52;
wire signed[31:0]    reg_activation_31_53;
wire signed[31:0]    reg_activation_31_54;
wire signed[31:0]    reg_activation_31_55;
wire signed[31:0]    reg_activation_31_56;
wire signed[31:0]    reg_activation_31_57;
wire signed[31:0]    reg_activation_31_58;
wire signed[31:0]    reg_activation_31_59;
wire signed[31:0]    reg_activation_31_60;
wire signed[31:0]    reg_activation_31_61;
wire signed[31:0]    reg_activation_31_62;
wire signed[31:0]    reg_activation_31_63;
wire signed[31:0]    reg_activation_32_0;
wire signed[31:0]    reg_activation_32_1;
wire signed[31:0]    reg_activation_32_2;
wire signed[31:0]    reg_activation_32_3;
wire signed[31:0]    reg_activation_32_4;
wire signed[31:0]    reg_activation_32_5;
wire signed[31:0]    reg_activation_32_6;
wire signed[31:0]    reg_activation_32_7;
wire signed[31:0]    reg_activation_32_8;
wire signed[31:0]    reg_activation_32_9;
wire signed[31:0]    reg_activation_32_10;
wire signed[31:0]    reg_activation_32_11;
wire signed[31:0]    reg_activation_32_12;
wire signed[31:0]    reg_activation_32_13;
wire signed[31:0]    reg_activation_32_14;
wire signed[31:0]    reg_activation_32_15;
wire signed[31:0]    reg_activation_32_16;
wire signed[31:0]    reg_activation_32_17;
wire signed[31:0]    reg_activation_32_18;
wire signed[31:0]    reg_activation_32_19;
wire signed[31:0]    reg_activation_32_20;
wire signed[31:0]    reg_activation_32_21;
wire signed[31:0]    reg_activation_32_22;
wire signed[31:0]    reg_activation_32_23;
wire signed[31:0]    reg_activation_32_24;
wire signed[31:0]    reg_activation_32_25;
wire signed[31:0]    reg_activation_32_26;
wire signed[31:0]    reg_activation_32_27;
wire signed[31:0]    reg_activation_32_28;
wire signed[31:0]    reg_activation_32_29;
wire signed[31:0]    reg_activation_32_30;
wire signed[31:0]    reg_activation_32_31;
wire signed[31:0]    reg_activation_32_32;
wire signed[31:0]    reg_activation_32_33;
wire signed[31:0]    reg_activation_32_34;
wire signed[31:0]    reg_activation_32_35;
wire signed[31:0]    reg_activation_32_36;
wire signed[31:0]    reg_activation_32_37;
wire signed[31:0]    reg_activation_32_38;
wire signed[31:0]    reg_activation_32_39;
wire signed[31:0]    reg_activation_32_40;
wire signed[31:0]    reg_activation_32_41;
wire signed[31:0]    reg_activation_32_42;
wire signed[31:0]    reg_activation_32_43;
wire signed[31:0]    reg_activation_32_44;
wire signed[31:0]    reg_activation_32_45;
wire signed[31:0]    reg_activation_32_46;
wire signed[31:0]    reg_activation_32_47;
wire signed[31:0]    reg_activation_32_48;
wire signed[31:0]    reg_activation_32_49;
wire signed[31:0]    reg_activation_32_50;
wire signed[31:0]    reg_activation_32_51;
wire signed[31:0]    reg_activation_32_52;
wire signed[31:0]    reg_activation_32_53;
wire signed[31:0]    reg_activation_32_54;
wire signed[31:0]    reg_activation_32_55;
wire signed[31:0]    reg_activation_32_56;
wire signed[31:0]    reg_activation_32_57;
wire signed[31:0]    reg_activation_32_58;
wire signed[31:0]    reg_activation_32_59;
wire signed[31:0]    reg_activation_32_60;
wire signed[31:0]    reg_activation_32_61;
wire signed[31:0]    reg_activation_32_62;
wire signed[31:0]    reg_activation_32_63;
wire signed[31:0]    reg_activation_33_0;
wire signed[31:0]    reg_activation_33_1;
wire signed[31:0]    reg_activation_33_2;
wire signed[31:0]    reg_activation_33_3;
wire signed[31:0]    reg_activation_33_4;
wire signed[31:0]    reg_activation_33_5;
wire signed[31:0]    reg_activation_33_6;
wire signed[31:0]    reg_activation_33_7;
wire signed[31:0]    reg_activation_33_8;
wire signed[31:0]    reg_activation_33_9;
wire signed[31:0]    reg_activation_33_10;
wire signed[31:0]    reg_activation_33_11;
wire signed[31:0]    reg_activation_33_12;
wire signed[31:0]    reg_activation_33_13;
wire signed[31:0]    reg_activation_33_14;
wire signed[31:0]    reg_activation_33_15;
wire signed[31:0]    reg_activation_33_16;
wire signed[31:0]    reg_activation_33_17;
wire signed[31:0]    reg_activation_33_18;
wire signed[31:0]    reg_activation_33_19;
wire signed[31:0]    reg_activation_33_20;
wire signed[31:0]    reg_activation_33_21;
wire signed[31:0]    reg_activation_33_22;
wire signed[31:0]    reg_activation_33_23;
wire signed[31:0]    reg_activation_33_24;
wire signed[31:0]    reg_activation_33_25;
wire signed[31:0]    reg_activation_33_26;
wire signed[31:0]    reg_activation_33_27;
wire signed[31:0]    reg_activation_33_28;
wire signed[31:0]    reg_activation_33_29;
wire signed[31:0]    reg_activation_33_30;
wire signed[31:0]    reg_activation_33_31;
wire signed[31:0]    reg_activation_33_32;
wire signed[31:0]    reg_activation_33_33;
wire signed[31:0]    reg_activation_33_34;
wire signed[31:0]    reg_activation_33_35;
wire signed[31:0]    reg_activation_33_36;
wire signed[31:0]    reg_activation_33_37;
wire signed[31:0]    reg_activation_33_38;
wire signed[31:0]    reg_activation_33_39;
wire signed[31:0]    reg_activation_33_40;
wire signed[31:0]    reg_activation_33_41;
wire signed[31:0]    reg_activation_33_42;
wire signed[31:0]    reg_activation_33_43;
wire signed[31:0]    reg_activation_33_44;
wire signed[31:0]    reg_activation_33_45;
wire signed[31:0]    reg_activation_33_46;
wire signed[31:0]    reg_activation_33_47;
wire signed[31:0]    reg_activation_33_48;
wire signed[31:0]    reg_activation_33_49;
wire signed[31:0]    reg_activation_33_50;
wire signed[31:0]    reg_activation_33_51;
wire signed[31:0]    reg_activation_33_52;
wire signed[31:0]    reg_activation_33_53;
wire signed[31:0]    reg_activation_33_54;
wire signed[31:0]    reg_activation_33_55;
wire signed[31:0]    reg_activation_33_56;
wire signed[31:0]    reg_activation_33_57;
wire signed[31:0]    reg_activation_33_58;
wire signed[31:0]    reg_activation_33_59;
wire signed[31:0]    reg_activation_33_60;
wire signed[31:0]    reg_activation_33_61;
wire signed[31:0]    reg_activation_33_62;
wire signed[31:0]    reg_activation_33_63;
wire signed[31:0]    reg_activation_34_0;
wire signed[31:0]    reg_activation_34_1;
wire signed[31:0]    reg_activation_34_2;
wire signed[31:0]    reg_activation_34_3;
wire signed[31:0]    reg_activation_34_4;
wire signed[31:0]    reg_activation_34_5;
wire signed[31:0]    reg_activation_34_6;
wire signed[31:0]    reg_activation_34_7;
wire signed[31:0]    reg_activation_34_8;
wire signed[31:0]    reg_activation_34_9;
wire signed[31:0]    reg_activation_34_10;
wire signed[31:0]    reg_activation_34_11;
wire signed[31:0]    reg_activation_34_12;
wire signed[31:0]    reg_activation_34_13;
wire signed[31:0]    reg_activation_34_14;
wire signed[31:0]    reg_activation_34_15;
wire signed[31:0]    reg_activation_34_16;
wire signed[31:0]    reg_activation_34_17;
wire signed[31:0]    reg_activation_34_18;
wire signed[31:0]    reg_activation_34_19;
wire signed[31:0]    reg_activation_34_20;
wire signed[31:0]    reg_activation_34_21;
wire signed[31:0]    reg_activation_34_22;
wire signed[31:0]    reg_activation_34_23;
wire signed[31:0]    reg_activation_34_24;
wire signed[31:0]    reg_activation_34_25;
wire signed[31:0]    reg_activation_34_26;
wire signed[31:0]    reg_activation_34_27;
wire signed[31:0]    reg_activation_34_28;
wire signed[31:0]    reg_activation_34_29;
wire signed[31:0]    reg_activation_34_30;
wire signed[31:0]    reg_activation_34_31;
wire signed[31:0]    reg_activation_34_32;
wire signed[31:0]    reg_activation_34_33;
wire signed[31:0]    reg_activation_34_34;
wire signed[31:0]    reg_activation_34_35;
wire signed[31:0]    reg_activation_34_36;
wire signed[31:0]    reg_activation_34_37;
wire signed[31:0]    reg_activation_34_38;
wire signed[31:0]    reg_activation_34_39;
wire signed[31:0]    reg_activation_34_40;
wire signed[31:0]    reg_activation_34_41;
wire signed[31:0]    reg_activation_34_42;
wire signed[31:0]    reg_activation_34_43;
wire signed[31:0]    reg_activation_34_44;
wire signed[31:0]    reg_activation_34_45;
wire signed[31:0]    reg_activation_34_46;
wire signed[31:0]    reg_activation_34_47;
wire signed[31:0]    reg_activation_34_48;
wire signed[31:0]    reg_activation_34_49;
wire signed[31:0]    reg_activation_34_50;
wire signed[31:0]    reg_activation_34_51;
wire signed[31:0]    reg_activation_34_52;
wire signed[31:0]    reg_activation_34_53;
wire signed[31:0]    reg_activation_34_54;
wire signed[31:0]    reg_activation_34_55;
wire signed[31:0]    reg_activation_34_56;
wire signed[31:0]    reg_activation_34_57;
wire signed[31:0]    reg_activation_34_58;
wire signed[31:0]    reg_activation_34_59;
wire signed[31:0]    reg_activation_34_60;
wire signed[31:0]    reg_activation_34_61;
wire signed[31:0]    reg_activation_34_62;
wire signed[31:0]    reg_activation_34_63;
wire signed[31:0]    reg_activation_35_0;
wire signed[31:0]    reg_activation_35_1;
wire signed[31:0]    reg_activation_35_2;
wire signed[31:0]    reg_activation_35_3;
wire signed[31:0]    reg_activation_35_4;
wire signed[31:0]    reg_activation_35_5;
wire signed[31:0]    reg_activation_35_6;
wire signed[31:0]    reg_activation_35_7;
wire signed[31:0]    reg_activation_35_8;
wire signed[31:0]    reg_activation_35_9;
wire signed[31:0]    reg_activation_35_10;
wire signed[31:0]    reg_activation_35_11;
wire signed[31:0]    reg_activation_35_12;
wire signed[31:0]    reg_activation_35_13;
wire signed[31:0]    reg_activation_35_14;
wire signed[31:0]    reg_activation_35_15;
wire signed[31:0]    reg_activation_35_16;
wire signed[31:0]    reg_activation_35_17;
wire signed[31:0]    reg_activation_35_18;
wire signed[31:0]    reg_activation_35_19;
wire signed[31:0]    reg_activation_35_20;
wire signed[31:0]    reg_activation_35_21;
wire signed[31:0]    reg_activation_35_22;
wire signed[31:0]    reg_activation_35_23;
wire signed[31:0]    reg_activation_35_24;
wire signed[31:0]    reg_activation_35_25;
wire signed[31:0]    reg_activation_35_26;
wire signed[31:0]    reg_activation_35_27;
wire signed[31:0]    reg_activation_35_28;
wire signed[31:0]    reg_activation_35_29;
wire signed[31:0]    reg_activation_35_30;
wire signed[31:0]    reg_activation_35_31;
wire signed[31:0]    reg_activation_35_32;
wire signed[31:0]    reg_activation_35_33;
wire signed[31:0]    reg_activation_35_34;
wire signed[31:0]    reg_activation_35_35;
wire signed[31:0]    reg_activation_35_36;
wire signed[31:0]    reg_activation_35_37;
wire signed[31:0]    reg_activation_35_38;
wire signed[31:0]    reg_activation_35_39;
wire signed[31:0]    reg_activation_35_40;
wire signed[31:0]    reg_activation_35_41;
wire signed[31:0]    reg_activation_35_42;
wire signed[31:0]    reg_activation_35_43;
wire signed[31:0]    reg_activation_35_44;
wire signed[31:0]    reg_activation_35_45;
wire signed[31:0]    reg_activation_35_46;
wire signed[31:0]    reg_activation_35_47;
wire signed[31:0]    reg_activation_35_48;
wire signed[31:0]    reg_activation_35_49;
wire signed[31:0]    reg_activation_35_50;
wire signed[31:0]    reg_activation_35_51;
wire signed[31:0]    reg_activation_35_52;
wire signed[31:0]    reg_activation_35_53;
wire signed[31:0]    reg_activation_35_54;
wire signed[31:0]    reg_activation_35_55;
wire signed[31:0]    reg_activation_35_56;
wire signed[31:0]    reg_activation_35_57;
wire signed[31:0]    reg_activation_35_58;
wire signed[31:0]    reg_activation_35_59;
wire signed[31:0]    reg_activation_35_60;
wire signed[31:0]    reg_activation_35_61;
wire signed[31:0]    reg_activation_35_62;
wire signed[31:0]    reg_activation_35_63;
wire signed[31:0]    reg_activation_36_0;
wire signed[31:0]    reg_activation_36_1;
wire signed[31:0]    reg_activation_36_2;
wire signed[31:0]    reg_activation_36_3;
wire signed[31:0]    reg_activation_36_4;
wire signed[31:0]    reg_activation_36_5;
wire signed[31:0]    reg_activation_36_6;
wire signed[31:0]    reg_activation_36_7;
wire signed[31:0]    reg_activation_36_8;
wire signed[31:0]    reg_activation_36_9;
wire signed[31:0]    reg_activation_36_10;
wire signed[31:0]    reg_activation_36_11;
wire signed[31:0]    reg_activation_36_12;
wire signed[31:0]    reg_activation_36_13;
wire signed[31:0]    reg_activation_36_14;
wire signed[31:0]    reg_activation_36_15;
wire signed[31:0]    reg_activation_36_16;
wire signed[31:0]    reg_activation_36_17;
wire signed[31:0]    reg_activation_36_18;
wire signed[31:0]    reg_activation_36_19;
wire signed[31:0]    reg_activation_36_20;
wire signed[31:0]    reg_activation_36_21;
wire signed[31:0]    reg_activation_36_22;
wire signed[31:0]    reg_activation_36_23;
wire signed[31:0]    reg_activation_36_24;
wire signed[31:0]    reg_activation_36_25;
wire signed[31:0]    reg_activation_36_26;
wire signed[31:0]    reg_activation_36_27;
wire signed[31:0]    reg_activation_36_28;
wire signed[31:0]    reg_activation_36_29;
wire signed[31:0]    reg_activation_36_30;
wire signed[31:0]    reg_activation_36_31;
wire signed[31:0]    reg_activation_36_32;
wire signed[31:0]    reg_activation_36_33;
wire signed[31:0]    reg_activation_36_34;
wire signed[31:0]    reg_activation_36_35;
wire signed[31:0]    reg_activation_36_36;
wire signed[31:0]    reg_activation_36_37;
wire signed[31:0]    reg_activation_36_38;
wire signed[31:0]    reg_activation_36_39;
wire signed[31:0]    reg_activation_36_40;
wire signed[31:0]    reg_activation_36_41;
wire signed[31:0]    reg_activation_36_42;
wire signed[31:0]    reg_activation_36_43;
wire signed[31:0]    reg_activation_36_44;
wire signed[31:0]    reg_activation_36_45;
wire signed[31:0]    reg_activation_36_46;
wire signed[31:0]    reg_activation_36_47;
wire signed[31:0]    reg_activation_36_48;
wire signed[31:0]    reg_activation_36_49;
wire signed[31:0]    reg_activation_36_50;
wire signed[31:0]    reg_activation_36_51;
wire signed[31:0]    reg_activation_36_52;
wire signed[31:0]    reg_activation_36_53;
wire signed[31:0]    reg_activation_36_54;
wire signed[31:0]    reg_activation_36_55;
wire signed[31:0]    reg_activation_36_56;
wire signed[31:0]    reg_activation_36_57;
wire signed[31:0]    reg_activation_36_58;
wire signed[31:0]    reg_activation_36_59;
wire signed[31:0]    reg_activation_36_60;
wire signed[31:0]    reg_activation_36_61;
wire signed[31:0]    reg_activation_36_62;
wire signed[31:0]    reg_activation_36_63;
wire signed[31:0]    reg_activation_37_0;
wire signed[31:0]    reg_activation_37_1;
wire signed[31:0]    reg_activation_37_2;
wire signed[31:0]    reg_activation_37_3;
wire signed[31:0]    reg_activation_37_4;
wire signed[31:0]    reg_activation_37_5;
wire signed[31:0]    reg_activation_37_6;
wire signed[31:0]    reg_activation_37_7;
wire signed[31:0]    reg_activation_37_8;
wire signed[31:0]    reg_activation_37_9;
wire signed[31:0]    reg_activation_37_10;
wire signed[31:0]    reg_activation_37_11;
wire signed[31:0]    reg_activation_37_12;
wire signed[31:0]    reg_activation_37_13;
wire signed[31:0]    reg_activation_37_14;
wire signed[31:0]    reg_activation_37_15;
wire signed[31:0]    reg_activation_37_16;
wire signed[31:0]    reg_activation_37_17;
wire signed[31:0]    reg_activation_37_18;
wire signed[31:0]    reg_activation_37_19;
wire signed[31:0]    reg_activation_37_20;
wire signed[31:0]    reg_activation_37_21;
wire signed[31:0]    reg_activation_37_22;
wire signed[31:0]    reg_activation_37_23;
wire signed[31:0]    reg_activation_37_24;
wire signed[31:0]    reg_activation_37_25;
wire signed[31:0]    reg_activation_37_26;
wire signed[31:0]    reg_activation_37_27;
wire signed[31:0]    reg_activation_37_28;
wire signed[31:0]    reg_activation_37_29;
wire signed[31:0]    reg_activation_37_30;
wire signed[31:0]    reg_activation_37_31;
wire signed[31:0]    reg_activation_37_32;
wire signed[31:0]    reg_activation_37_33;
wire signed[31:0]    reg_activation_37_34;
wire signed[31:0]    reg_activation_37_35;
wire signed[31:0]    reg_activation_37_36;
wire signed[31:0]    reg_activation_37_37;
wire signed[31:0]    reg_activation_37_38;
wire signed[31:0]    reg_activation_37_39;
wire signed[31:0]    reg_activation_37_40;
wire signed[31:0]    reg_activation_37_41;
wire signed[31:0]    reg_activation_37_42;
wire signed[31:0]    reg_activation_37_43;
wire signed[31:0]    reg_activation_37_44;
wire signed[31:0]    reg_activation_37_45;
wire signed[31:0]    reg_activation_37_46;
wire signed[31:0]    reg_activation_37_47;
wire signed[31:0]    reg_activation_37_48;
wire signed[31:0]    reg_activation_37_49;
wire signed[31:0]    reg_activation_37_50;
wire signed[31:0]    reg_activation_37_51;
wire signed[31:0]    reg_activation_37_52;
wire signed[31:0]    reg_activation_37_53;
wire signed[31:0]    reg_activation_37_54;
wire signed[31:0]    reg_activation_37_55;
wire signed[31:0]    reg_activation_37_56;
wire signed[31:0]    reg_activation_37_57;
wire signed[31:0]    reg_activation_37_58;
wire signed[31:0]    reg_activation_37_59;
wire signed[31:0]    reg_activation_37_60;
wire signed[31:0]    reg_activation_37_61;
wire signed[31:0]    reg_activation_37_62;
wire signed[31:0]    reg_activation_37_63;
wire signed[31:0]    reg_activation_38_0;
wire signed[31:0]    reg_activation_38_1;
wire signed[31:0]    reg_activation_38_2;
wire signed[31:0]    reg_activation_38_3;
wire signed[31:0]    reg_activation_38_4;
wire signed[31:0]    reg_activation_38_5;
wire signed[31:0]    reg_activation_38_6;
wire signed[31:0]    reg_activation_38_7;
wire signed[31:0]    reg_activation_38_8;
wire signed[31:0]    reg_activation_38_9;
wire signed[31:0]    reg_activation_38_10;
wire signed[31:0]    reg_activation_38_11;
wire signed[31:0]    reg_activation_38_12;
wire signed[31:0]    reg_activation_38_13;
wire signed[31:0]    reg_activation_38_14;
wire signed[31:0]    reg_activation_38_15;
wire signed[31:0]    reg_activation_38_16;
wire signed[31:0]    reg_activation_38_17;
wire signed[31:0]    reg_activation_38_18;
wire signed[31:0]    reg_activation_38_19;
wire signed[31:0]    reg_activation_38_20;
wire signed[31:0]    reg_activation_38_21;
wire signed[31:0]    reg_activation_38_22;
wire signed[31:0]    reg_activation_38_23;
wire signed[31:0]    reg_activation_38_24;
wire signed[31:0]    reg_activation_38_25;
wire signed[31:0]    reg_activation_38_26;
wire signed[31:0]    reg_activation_38_27;
wire signed[31:0]    reg_activation_38_28;
wire signed[31:0]    reg_activation_38_29;
wire signed[31:0]    reg_activation_38_30;
wire signed[31:0]    reg_activation_38_31;
wire signed[31:0]    reg_activation_38_32;
wire signed[31:0]    reg_activation_38_33;
wire signed[31:0]    reg_activation_38_34;
wire signed[31:0]    reg_activation_38_35;
wire signed[31:0]    reg_activation_38_36;
wire signed[31:0]    reg_activation_38_37;
wire signed[31:0]    reg_activation_38_38;
wire signed[31:0]    reg_activation_38_39;
wire signed[31:0]    reg_activation_38_40;
wire signed[31:0]    reg_activation_38_41;
wire signed[31:0]    reg_activation_38_42;
wire signed[31:0]    reg_activation_38_43;
wire signed[31:0]    reg_activation_38_44;
wire signed[31:0]    reg_activation_38_45;
wire signed[31:0]    reg_activation_38_46;
wire signed[31:0]    reg_activation_38_47;
wire signed[31:0]    reg_activation_38_48;
wire signed[31:0]    reg_activation_38_49;
wire signed[31:0]    reg_activation_38_50;
wire signed[31:0]    reg_activation_38_51;
wire signed[31:0]    reg_activation_38_52;
wire signed[31:0]    reg_activation_38_53;
wire signed[31:0]    reg_activation_38_54;
wire signed[31:0]    reg_activation_38_55;
wire signed[31:0]    reg_activation_38_56;
wire signed[31:0]    reg_activation_38_57;
wire signed[31:0]    reg_activation_38_58;
wire signed[31:0]    reg_activation_38_59;
wire signed[31:0]    reg_activation_38_60;
wire signed[31:0]    reg_activation_38_61;
wire signed[31:0]    reg_activation_38_62;
wire signed[31:0]    reg_activation_38_63;
wire signed[31:0]    reg_activation_39_0;
wire signed[31:0]    reg_activation_39_1;
wire signed[31:0]    reg_activation_39_2;
wire signed[31:0]    reg_activation_39_3;
wire signed[31:0]    reg_activation_39_4;
wire signed[31:0]    reg_activation_39_5;
wire signed[31:0]    reg_activation_39_6;
wire signed[31:0]    reg_activation_39_7;
wire signed[31:0]    reg_activation_39_8;
wire signed[31:0]    reg_activation_39_9;
wire signed[31:0]    reg_activation_39_10;
wire signed[31:0]    reg_activation_39_11;
wire signed[31:0]    reg_activation_39_12;
wire signed[31:0]    reg_activation_39_13;
wire signed[31:0]    reg_activation_39_14;
wire signed[31:0]    reg_activation_39_15;
wire signed[31:0]    reg_activation_39_16;
wire signed[31:0]    reg_activation_39_17;
wire signed[31:0]    reg_activation_39_18;
wire signed[31:0]    reg_activation_39_19;
wire signed[31:0]    reg_activation_39_20;
wire signed[31:0]    reg_activation_39_21;
wire signed[31:0]    reg_activation_39_22;
wire signed[31:0]    reg_activation_39_23;
wire signed[31:0]    reg_activation_39_24;
wire signed[31:0]    reg_activation_39_25;
wire signed[31:0]    reg_activation_39_26;
wire signed[31:0]    reg_activation_39_27;
wire signed[31:0]    reg_activation_39_28;
wire signed[31:0]    reg_activation_39_29;
wire signed[31:0]    reg_activation_39_30;
wire signed[31:0]    reg_activation_39_31;
wire signed[31:0]    reg_activation_39_32;
wire signed[31:0]    reg_activation_39_33;
wire signed[31:0]    reg_activation_39_34;
wire signed[31:0]    reg_activation_39_35;
wire signed[31:0]    reg_activation_39_36;
wire signed[31:0]    reg_activation_39_37;
wire signed[31:0]    reg_activation_39_38;
wire signed[31:0]    reg_activation_39_39;
wire signed[31:0]    reg_activation_39_40;
wire signed[31:0]    reg_activation_39_41;
wire signed[31:0]    reg_activation_39_42;
wire signed[31:0]    reg_activation_39_43;
wire signed[31:0]    reg_activation_39_44;
wire signed[31:0]    reg_activation_39_45;
wire signed[31:0]    reg_activation_39_46;
wire signed[31:0]    reg_activation_39_47;
wire signed[31:0]    reg_activation_39_48;
wire signed[31:0]    reg_activation_39_49;
wire signed[31:0]    reg_activation_39_50;
wire signed[31:0]    reg_activation_39_51;
wire signed[31:0]    reg_activation_39_52;
wire signed[31:0]    reg_activation_39_53;
wire signed[31:0]    reg_activation_39_54;
wire signed[31:0]    reg_activation_39_55;
wire signed[31:0]    reg_activation_39_56;
wire signed[31:0]    reg_activation_39_57;
wire signed[31:0]    reg_activation_39_58;
wire signed[31:0]    reg_activation_39_59;
wire signed[31:0]    reg_activation_39_60;
wire signed[31:0]    reg_activation_39_61;
wire signed[31:0]    reg_activation_39_62;
wire signed[31:0]    reg_activation_39_63;
wire signed[31:0]    reg_activation_40_0;
wire signed[31:0]    reg_activation_40_1;
wire signed[31:0]    reg_activation_40_2;
wire signed[31:0]    reg_activation_40_3;
wire signed[31:0]    reg_activation_40_4;
wire signed[31:0]    reg_activation_40_5;
wire signed[31:0]    reg_activation_40_6;
wire signed[31:0]    reg_activation_40_7;
wire signed[31:0]    reg_activation_40_8;
wire signed[31:0]    reg_activation_40_9;
wire signed[31:0]    reg_activation_40_10;
wire signed[31:0]    reg_activation_40_11;
wire signed[31:0]    reg_activation_40_12;
wire signed[31:0]    reg_activation_40_13;
wire signed[31:0]    reg_activation_40_14;
wire signed[31:0]    reg_activation_40_15;
wire signed[31:0]    reg_activation_40_16;
wire signed[31:0]    reg_activation_40_17;
wire signed[31:0]    reg_activation_40_18;
wire signed[31:0]    reg_activation_40_19;
wire signed[31:0]    reg_activation_40_20;
wire signed[31:0]    reg_activation_40_21;
wire signed[31:0]    reg_activation_40_22;
wire signed[31:0]    reg_activation_40_23;
wire signed[31:0]    reg_activation_40_24;
wire signed[31:0]    reg_activation_40_25;
wire signed[31:0]    reg_activation_40_26;
wire signed[31:0]    reg_activation_40_27;
wire signed[31:0]    reg_activation_40_28;
wire signed[31:0]    reg_activation_40_29;
wire signed[31:0]    reg_activation_40_30;
wire signed[31:0]    reg_activation_40_31;
wire signed[31:0]    reg_activation_40_32;
wire signed[31:0]    reg_activation_40_33;
wire signed[31:0]    reg_activation_40_34;
wire signed[31:0]    reg_activation_40_35;
wire signed[31:0]    reg_activation_40_36;
wire signed[31:0]    reg_activation_40_37;
wire signed[31:0]    reg_activation_40_38;
wire signed[31:0]    reg_activation_40_39;
wire signed[31:0]    reg_activation_40_40;
wire signed[31:0]    reg_activation_40_41;
wire signed[31:0]    reg_activation_40_42;
wire signed[31:0]    reg_activation_40_43;
wire signed[31:0]    reg_activation_40_44;
wire signed[31:0]    reg_activation_40_45;
wire signed[31:0]    reg_activation_40_46;
wire signed[31:0]    reg_activation_40_47;
wire signed[31:0]    reg_activation_40_48;
wire signed[31:0]    reg_activation_40_49;
wire signed[31:0]    reg_activation_40_50;
wire signed[31:0]    reg_activation_40_51;
wire signed[31:0]    reg_activation_40_52;
wire signed[31:0]    reg_activation_40_53;
wire signed[31:0]    reg_activation_40_54;
wire signed[31:0]    reg_activation_40_55;
wire signed[31:0]    reg_activation_40_56;
wire signed[31:0]    reg_activation_40_57;
wire signed[31:0]    reg_activation_40_58;
wire signed[31:0]    reg_activation_40_59;
wire signed[31:0]    reg_activation_40_60;
wire signed[31:0]    reg_activation_40_61;
wire signed[31:0]    reg_activation_40_62;
wire signed[31:0]    reg_activation_40_63;
wire signed[31:0]    reg_activation_41_0;
wire signed[31:0]    reg_activation_41_1;
wire signed[31:0]    reg_activation_41_2;
wire signed[31:0]    reg_activation_41_3;
wire signed[31:0]    reg_activation_41_4;
wire signed[31:0]    reg_activation_41_5;
wire signed[31:0]    reg_activation_41_6;
wire signed[31:0]    reg_activation_41_7;
wire signed[31:0]    reg_activation_41_8;
wire signed[31:0]    reg_activation_41_9;
wire signed[31:0]    reg_activation_41_10;
wire signed[31:0]    reg_activation_41_11;
wire signed[31:0]    reg_activation_41_12;
wire signed[31:0]    reg_activation_41_13;
wire signed[31:0]    reg_activation_41_14;
wire signed[31:0]    reg_activation_41_15;
wire signed[31:0]    reg_activation_41_16;
wire signed[31:0]    reg_activation_41_17;
wire signed[31:0]    reg_activation_41_18;
wire signed[31:0]    reg_activation_41_19;
wire signed[31:0]    reg_activation_41_20;
wire signed[31:0]    reg_activation_41_21;
wire signed[31:0]    reg_activation_41_22;
wire signed[31:0]    reg_activation_41_23;
wire signed[31:0]    reg_activation_41_24;
wire signed[31:0]    reg_activation_41_25;
wire signed[31:0]    reg_activation_41_26;
wire signed[31:0]    reg_activation_41_27;
wire signed[31:0]    reg_activation_41_28;
wire signed[31:0]    reg_activation_41_29;
wire signed[31:0]    reg_activation_41_30;
wire signed[31:0]    reg_activation_41_31;
wire signed[31:0]    reg_activation_41_32;
wire signed[31:0]    reg_activation_41_33;
wire signed[31:0]    reg_activation_41_34;
wire signed[31:0]    reg_activation_41_35;
wire signed[31:0]    reg_activation_41_36;
wire signed[31:0]    reg_activation_41_37;
wire signed[31:0]    reg_activation_41_38;
wire signed[31:0]    reg_activation_41_39;
wire signed[31:0]    reg_activation_41_40;
wire signed[31:0]    reg_activation_41_41;
wire signed[31:0]    reg_activation_41_42;
wire signed[31:0]    reg_activation_41_43;
wire signed[31:0]    reg_activation_41_44;
wire signed[31:0]    reg_activation_41_45;
wire signed[31:0]    reg_activation_41_46;
wire signed[31:0]    reg_activation_41_47;
wire signed[31:0]    reg_activation_41_48;
wire signed[31:0]    reg_activation_41_49;
wire signed[31:0]    reg_activation_41_50;
wire signed[31:0]    reg_activation_41_51;
wire signed[31:0]    reg_activation_41_52;
wire signed[31:0]    reg_activation_41_53;
wire signed[31:0]    reg_activation_41_54;
wire signed[31:0]    reg_activation_41_55;
wire signed[31:0]    reg_activation_41_56;
wire signed[31:0]    reg_activation_41_57;
wire signed[31:0]    reg_activation_41_58;
wire signed[31:0]    reg_activation_41_59;
wire signed[31:0]    reg_activation_41_60;
wire signed[31:0]    reg_activation_41_61;
wire signed[31:0]    reg_activation_41_62;
wire signed[31:0]    reg_activation_41_63;
wire signed[31:0]    reg_activation_42_0;
wire signed[31:0]    reg_activation_42_1;
wire signed[31:0]    reg_activation_42_2;
wire signed[31:0]    reg_activation_42_3;
wire signed[31:0]    reg_activation_42_4;
wire signed[31:0]    reg_activation_42_5;
wire signed[31:0]    reg_activation_42_6;
wire signed[31:0]    reg_activation_42_7;
wire signed[31:0]    reg_activation_42_8;
wire signed[31:0]    reg_activation_42_9;
wire signed[31:0]    reg_activation_42_10;
wire signed[31:0]    reg_activation_42_11;
wire signed[31:0]    reg_activation_42_12;
wire signed[31:0]    reg_activation_42_13;
wire signed[31:0]    reg_activation_42_14;
wire signed[31:0]    reg_activation_42_15;
wire signed[31:0]    reg_activation_42_16;
wire signed[31:0]    reg_activation_42_17;
wire signed[31:0]    reg_activation_42_18;
wire signed[31:0]    reg_activation_42_19;
wire signed[31:0]    reg_activation_42_20;
wire signed[31:0]    reg_activation_42_21;
wire signed[31:0]    reg_activation_42_22;
wire signed[31:0]    reg_activation_42_23;
wire signed[31:0]    reg_activation_42_24;
wire signed[31:0]    reg_activation_42_25;
wire signed[31:0]    reg_activation_42_26;
wire signed[31:0]    reg_activation_42_27;
wire signed[31:0]    reg_activation_42_28;
wire signed[31:0]    reg_activation_42_29;
wire signed[31:0]    reg_activation_42_30;
wire signed[31:0]    reg_activation_42_31;
wire signed[31:0]    reg_activation_42_32;
wire signed[31:0]    reg_activation_42_33;
wire signed[31:0]    reg_activation_42_34;
wire signed[31:0]    reg_activation_42_35;
wire signed[31:0]    reg_activation_42_36;
wire signed[31:0]    reg_activation_42_37;
wire signed[31:0]    reg_activation_42_38;
wire signed[31:0]    reg_activation_42_39;
wire signed[31:0]    reg_activation_42_40;
wire signed[31:0]    reg_activation_42_41;
wire signed[31:0]    reg_activation_42_42;
wire signed[31:0]    reg_activation_42_43;
wire signed[31:0]    reg_activation_42_44;
wire signed[31:0]    reg_activation_42_45;
wire signed[31:0]    reg_activation_42_46;
wire signed[31:0]    reg_activation_42_47;
wire signed[31:0]    reg_activation_42_48;
wire signed[31:0]    reg_activation_42_49;
wire signed[31:0]    reg_activation_42_50;
wire signed[31:0]    reg_activation_42_51;
wire signed[31:0]    reg_activation_42_52;
wire signed[31:0]    reg_activation_42_53;
wire signed[31:0]    reg_activation_42_54;
wire signed[31:0]    reg_activation_42_55;
wire signed[31:0]    reg_activation_42_56;
wire signed[31:0]    reg_activation_42_57;
wire signed[31:0]    reg_activation_42_58;
wire signed[31:0]    reg_activation_42_59;
wire signed[31:0]    reg_activation_42_60;
wire signed[31:0]    reg_activation_42_61;
wire signed[31:0]    reg_activation_42_62;
wire signed[31:0]    reg_activation_42_63;
wire signed[31:0]    reg_activation_43_0;
wire signed[31:0]    reg_activation_43_1;
wire signed[31:0]    reg_activation_43_2;
wire signed[31:0]    reg_activation_43_3;
wire signed[31:0]    reg_activation_43_4;
wire signed[31:0]    reg_activation_43_5;
wire signed[31:0]    reg_activation_43_6;
wire signed[31:0]    reg_activation_43_7;
wire signed[31:0]    reg_activation_43_8;
wire signed[31:0]    reg_activation_43_9;
wire signed[31:0]    reg_activation_43_10;
wire signed[31:0]    reg_activation_43_11;
wire signed[31:0]    reg_activation_43_12;
wire signed[31:0]    reg_activation_43_13;
wire signed[31:0]    reg_activation_43_14;
wire signed[31:0]    reg_activation_43_15;
wire signed[31:0]    reg_activation_43_16;
wire signed[31:0]    reg_activation_43_17;
wire signed[31:0]    reg_activation_43_18;
wire signed[31:0]    reg_activation_43_19;
wire signed[31:0]    reg_activation_43_20;
wire signed[31:0]    reg_activation_43_21;
wire signed[31:0]    reg_activation_43_22;
wire signed[31:0]    reg_activation_43_23;
wire signed[31:0]    reg_activation_43_24;
wire signed[31:0]    reg_activation_43_25;
wire signed[31:0]    reg_activation_43_26;
wire signed[31:0]    reg_activation_43_27;
wire signed[31:0]    reg_activation_43_28;
wire signed[31:0]    reg_activation_43_29;
wire signed[31:0]    reg_activation_43_30;
wire signed[31:0]    reg_activation_43_31;
wire signed[31:0]    reg_activation_43_32;
wire signed[31:0]    reg_activation_43_33;
wire signed[31:0]    reg_activation_43_34;
wire signed[31:0]    reg_activation_43_35;
wire signed[31:0]    reg_activation_43_36;
wire signed[31:0]    reg_activation_43_37;
wire signed[31:0]    reg_activation_43_38;
wire signed[31:0]    reg_activation_43_39;
wire signed[31:0]    reg_activation_43_40;
wire signed[31:0]    reg_activation_43_41;
wire signed[31:0]    reg_activation_43_42;
wire signed[31:0]    reg_activation_43_43;
wire signed[31:0]    reg_activation_43_44;
wire signed[31:0]    reg_activation_43_45;
wire signed[31:0]    reg_activation_43_46;
wire signed[31:0]    reg_activation_43_47;
wire signed[31:0]    reg_activation_43_48;
wire signed[31:0]    reg_activation_43_49;
wire signed[31:0]    reg_activation_43_50;
wire signed[31:0]    reg_activation_43_51;
wire signed[31:0]    reg_activation_43_52;
wire signed[31:0]    reg_activation_43_53;
wire signed[31:0]    reg_activation_43_54;
wire signed[31:0]    reg_activation_43_55;
wire signed[31:0]    reg_activation_43_56;
wire signed[31:0]    reg_activation_43_57;
wire signed[31:0]    reg_activation_43_58;
wire signed[31:0]    reg_activation_43_59;
wire signed[31:0]    reg_activation_43_60;
wire signed[31:0]    reg_activation_43_61;
wire signed[31:0]    reg_activation_43_62;
wire signed[31:0]    reg_activation_43_63;
wire signed[31:0]    reg_activation_44_0;
wire signed[31:0]    reg_activation_44_1;
wire signed[31:0]    reg_activation_44_2;
wire signed[31:0]    reg_activation_44_3;
wire signed[31:0]    reg_activation_44_4;
wire signed[31:0]    reg_activation_44_5;
wire signed[31:0]    reg_activation_44_6;
wire signed[31:0]    reg_activation_44_7;
wire signed[31:0]    reg_activation_44_8;
wire signed[31:0]    reg_activation_44_9;
wire signed[31:0]    reg_activation_44_10;
wire signed[31:0]    reg_activation_44_11;
wire signed[31:0]    reg_activation_44_12;
wire signed[31:0]    reg_activation_44_13;
wire signed[31:0]    reg_activation_44_14;
wire signed[31:0]    reg_activation_44_15;
wire signed[31:0]    reg_activation_44_16;
wire signed[31:0]    reg_activation_44_17;
wire signed[31:0]    reg_activation_44_18;
wire signed[31:0]    reg_activation_44_19;
wire signed[31:0]    reg_activation_44_20;
wire signed[31:0]    reg_activation_44_21;
wire signed[31:0]    reg_activation_44_22;
wire signed[31:0]    reg_activation_44_23;
wire signed[31:0]    reg_activation_44_24;
wire signed[31:0]    reg_activation_44_25;
wire signed[31:0]    reg_activation_44_26;
wire signed[31:0]    reg_activation_44_27;
wire signed[31:0]    reg_activation_44_28;
wire signed[31:0]    reg_activation_44_29;
wire signed[31:0]    reg_activation_44_30;
wire signed[31:0]    reg_activation_44_31;
wire signed[31:0]    reg_activation_44_32;
wire signed[31:0]    reg_activation_44_33;
wire signed[31:0]    reg_activation_44_34;
wire signed[31:0]    reg_activation_44_35;
wire signed[31:0]    reg_activation_44_36;
wire signed[31:0]    reg_activation_44_37;
wire signed[31:0]    reg_activation_44_38;
wire signed[31:0]    reg_activation_44_39;
wire signed[31:0]    reg_activation_44_40;
wire signed[31:0]    reg_activation_44_41;
wire signed[31:0]    reg_activation_44_42;
wire signed[31:0]    reg_activation_44_43;
wire signed[31:0]    reg_activation_44_44;
wire signed[31:0]    reg_activation_44_45;
wire signed[31:0]    reg_activation_44_46;
wire signed[31:0]    reg_activation_44_47;
wire signed[31:0]    reg_activation_44_48;
wire signed[31:0]    reg_activation_44_49;
wire signed[31:0]    reg_activation_44_50;
wire signed[31:0]    reg_activation_44_51;
wire signed[31:0]    reg_activation_44_52;
wire signed[31:0]    reg_activation_44_53;
wire signed[31:0]    reg_activation_44_54;
wire signed[31:0]    reg_activation_44_55;
wire signed[31:0]    reg_activation_44_56;
wire signed[31:0]    reg_activation_44_57;
wire signed[31:0]    reg_activation_44_58;
wire signed[31:0]    reg_activation_44_59;
wire signed[31:0]    reg_activation_44_60;
wire signed[31:0]    reg_activation_44_61;
wire signed[31:0]    reg_activation_44_62;
wire signed[31:0]    reg_activation_44_63;
wire signed[31:0]    reg_activation_45_0;
wire signed[31:0]    reg_activation_45_1;
wire signed[31:0]    reg_activation_45_2;
wire signed[31:0]    reg_activation_45_3;
wire signed[31:0]    reg_activation_45_4;
wire signed[31:0]    reg_activation_45_5;
wire signed[31:0]    reg_activation_45_6;
wire signed[31:0]    reg_activation_45_7;
wire signed[31:0]    reg_activation_45_8;
wire signed[31:0]    reg_activation_45_9;
wire signed[31:0]    reg_activation_45_10;
wire signed[31:0]    reg_activation_45_11;
wire signed[31:0]    reg_activation_45_12;
wire signed[31:0]    reg_activation_45_13;
wire signed[31:0]    reg_activation_45_14;
wire signed[31:0]    reg_activation_45_15;
wire signed[31:0]    reg_activation_45_16;
wire signed[31:0]    reg_activation_45_17;
wire signed[31:0]    reg_activation_45_18;
wire signed[31:0]    reg_activation_45_19;
wire signed[31:0]    reg_activation_45_20;
wire signed[31:0]    reg_activation_45_21;
wire signed[31:0]    reg_activation_45_22;
wire signed[31:0]    reg_activation_45_23;
wire signed[31:0]    reg_activation_45_24;
wire signed[31:0]    reg_activation_45_25;
wire signed[31:0]    reg_activation_45_26;
wire signed[31:0]    reg_activation_45_27;
wire signed[31:0]    reg_activation_45_28;
wire signed[31:0]    reg_activation_45_29;
wire signed[31:0]    reg_activation_45_30;
wire signed[31:0]    reg_activation_45_31;
wire signed[31:0]    reg_activation_45_32;
wire signed[31:0]    reg_activation_45_33;
wire signed[31:0]    reg_activation_45_34;
wire signed[31:0]    reg_activation_45_35;
wire signed[31:0]    reg_activation_45_36;
wire signed[31:0]    reg_activation_45_37;
wire signed[31:0]    reg_activation_45_38;
wire signed[31:0]    reg_activation_45_39;
wire signed[31:0]    reg_activation_45_40;
wire signed[31:0]    reg_activation_45_41;
wire signed[31:0]    reg_activation_45_42;
wire signed[31:0]    reg_activation_45_43;
wire signed[31:0]    reg_activation_45_44;
wire signed[31:0]    reg_activation_45_45;
wire signed[31:0]    reg_activation_45_46;
wire signed[31:0]    reg_activation_45_47;
wire signed[31:0]    reg_activation_45_48;
wire signed[31:0]    reg_activation_45_49;
wire signed[31:0]    reg_activation_45_50;
wire signed[31:0]    reg_activation_45_51;
wire signed[31:0]    reg_activation_45_52;
wire signed[31:0]    reg_activation_45_53;
wire signed[31:0]    reg_activation_45_54;
wire signed[31:0]    reg_activation_45_55;
wire signed[31:0]    reg_activation_45_56;
wire signed[31:0]    reg_activation_45_57;
wire signed[31:0]    reg_activation_45_58;
wire signed[31:0]    reg_activation_45_59;
wire signed[31:0]    reg_activation_45_60;
wire signed[31:0]    reg_activation_45_61;
wire signed[31:0]    reg_activation_45_62;
wire signed[31:0]    reg_activation_45_63;
wire signed[31:0]    reg_activation_46_0;
wire signed[31:0]    reg_activation_46_1;
wire signed[31:0]    reg_activation_46_2;
wire signed[31:0]    reg_activation_46_3;
wire signed[31:0]    reg_activation_46_4;
wire signed[31:0]    reg_activation_46_5;
wire signed[31:0]    reg_activation_46_6;
wire signed[31:0]    reg_activation_46_7;
wire signed[31:0]    reg_activation_46_8;
wire signed[31:0]    reg_activation_46_9;
wire signed[31:0]    reg_activation_46_10;
wire signed[31:0]    reg_activation_46_11;
wire signed[31:0]    reg_activation_46_12;
wire signed[31:0]    reg_activation_46_13;
wire signed[31:0]    reg_activation_46_14;
wire signed[31:0]    reg_activation_46_15;
wire signed[31:0]    reg_activation_46_16;
wire signed[31:0]    reg_activation_46_17;
wire signed[31:0]    reg_activation_46_18;
wire signed[31:0]    reg_activation_46_19;
wire signed[31:0]    reg_activation_46_20;
wire signed[31:0]    reg_activation_46_21;
wire signed[31:0]    reg_activation_46_22;
wire signed[31:0]    reg_activation_46_23;
wire signed[31:0]    reg_activation_46_24;
wire signed[31:0]    reg_activation_46_25;
wire signed[31:0]    reg_activation_46_26;
wire signed[31:0]    reg_activation_46_27;
wire signed[31:0]    reg_activation_46_28;
wire signed[31:0]    reg_activation_46_29;
wire signed[31:0]    reg_activation_46_30;
wire signed[31:0]    reg_activation_46_31;
wire signed[31:0]    reg_activation_46_32;
wire signed[31:0]    reg_activation_46_33;
wire signed[31:0]    reg_activation_46_34;
wire signed[31:0]    reg_activation_46_35;
wire signed[31:0]    reg_activation_46_36;
wire signed[31:0]    reg_activation_46_37;
wire signed[31:0]    reg_activation_46_38;
wire signed[31:0]    reg_activation_46_39;
wire signed[31:0]    reg_activation_46_40;
wire signed[31:0]    reg_activation_46_41;
wire signed[31:0]    reg_activation_46_42;
wire signed[31:0]    reg_activation_46_43;
wire signed[31:0]    reg_activation_46_44;
wire signed[31:0]    reg_activation_46_45;
wire signed[31:0]    reg_activation_46_46;
wire signed[31:0]    reg_activation_46_47;
wire signed[31:0]    reg_activation_46_48;
wire signed[31:0]    reg_activation_46_49;
wire signed[31:0]    reg_activation_46_50;
wire signed[31:0]    reg_activation_46_51;
wire signed[31:0]    reg_activation_46_52;
wire signed[31:0]    reg_activation_46_53;
wire signed[31:0]    reg_activation_46_54;
wire signed[31:0]    reg_activation_46_55;
wire signed[31:0]    reg_activation_46_56;
wire signed[31:0]    reg_activation_46_57;
wire signed[31:0]    reg_activation_46_58;
wire signed[31:0]    reg_activation_46_59;
wire signed[31:0]    reg_activation_46_60;
wire signed[31:0]    reg_activation_46_61;
wire signed[31:0]    reg_activation_46_62;
wire signed[31:0]    reg_activation_46_63;
wire signed[31:0]    reg_activation_47_0;
wire signed[31:0]    reg_activation_47_1;
wire signed[31:0]    reg_activation_47_2;
wire signed[31:0]    reg_activation_47_3;
wire signed[31:0]    reg_activation_47_4;
wire signed[31:0]    reg_activation_47_5;
wire signed[31:0]    reg_activation_47_6;
wire signed[31:0]    reg_activation_47_7;
wire signed[31:0]    reg_activation_47_8;
wire signed[31:0]    reg_activation_47_9;
wire signed[31:0]    reg_activation_47_10;
wire signed[31:0]    reg_activation_47_11;
wire signed[31:0]    reg_activation_47_12;
wire signed[31:0]    reg_activation_47_13;
wire signed[31:0]    reg_activation_47_14;
wire signed[31:0]    reg_activation_47_15;
wire signed[31:0]    reg_activation_47_16;
wire signed[31:0]    reg_activation_47_17;
wire signed[31:0]    reg_activation_47_18;
wire signed[31:0]    reg_activation_47_19;
wire signed[31:0]    reg_activation_47_20;
wire signed[31:0]    reg_activation_47_21;
wire signed[31:0]    reg_activation_47_22;
wire signed[31:0]    reg_activation_47_23;
wire signed[31:0]    reg_activation_47_24;
wire signed[31:0]    reg_activation_47_25;
wire signed[31:0]    reg_activation_47_26;
wire signed[31:0]    reg_activation_47_27;
wire signed[31:0]    reg_activation_47_28;
wire signed[31:0]    reg_activation_47_29;
wire signed[31:0]    reg_activation_47_30;
wire signed[31:0]    reg_activation_47_31;
wire signed[31:0]    reg_activation_47_32;
wire signed[31:0]    reg_activation_47_33;
wire signed[31:0]    reg_activation_47_34;
wire signed[31:0]    reg_activation_47_35;
wire signed[31:0]    reg_activation_47_36;
wire signed[31:0]    reg_activation_47_37;
wire signed[31:0]    reg_activation_47_38;
wire signed[31:0]    reg_activation_47_39;
wire signed[31:0]    reg_activation_47_40;
wire signed[31:0]    reg_activation_47_41;
wire signed[31:0]    reg_activation_47_42;
wire signed[31:0]    reg_activation_47_43;
wire signed[31:0]    reg_activation_47_44;
wire signed[31:0]    reg_activation_47_45;
wire signed[31:0]    reg_activation_47_46;
wire signed[31:0]    reg_activation_47_47;
wire signed[31:0]    reg_activation_47_48;
wire signed[31:0]    reg_activation_47_49;
wire signed[31:0]    reg_activation_47_50;
wire signed[31:0]    reg_activation_47_51;
wire signed[31:0]    reg_activation_47_52;
wire signed[31:0]    reg_activation_47_53;
wire signed[31:0]    reg_activation_47_54;
wire signed[31:0]    reg_activation_47_55;
wire signed[31:0]    reg_activation_47_56;
wire signed[31:0]    reg_activation_47_57;
wire signed[31:0]    reg_activation_47_58;
wire signed[31:0]    reg_activation_47_59;
wire signed[31:0]    reg_activation_47_60;
wire signed[31:0]    reg_activation_47_61;
wire signed[31:0]    reg_activation_47_62;
wire signed[31:0]    reg_activation_47_63;
wire signed[31:0]    reg_activation_48_0;
wire signed[31:0]    reg_activation_48_1;
wire signed[31:0]    reg_activation_48_2;
wire signed[31:0]    reg_activation_48_3;
wire signed[31:0]    reg_activation_48_4;
wire signed[31:0]    reg_activation_48_5;
wire signed[31:0]    reg_activation_48_6;
wire signed[31:0]    reg_activation_48_7;
wire signed[31:0]    reg_activation_48_8;
wire signed[31:0]    reg_activation_48_9;
wire signed[31:0]    reg_activation_48_10;
wire signed[31:0]    reg_activation_48_11;
wire signed[31:0]    reg_activation_48_12;
wire signed[31:0]    reg_activation_48_13;
wire signed[31:0]    reg_activation_48_14;
wire signed[31:0]    reg_activation_48_15;
wire signed[31:0]    reg_activation_48_16;
wire signed[31:0]    reg_activation_48_17;
wire signed[31:0]    reg_activation_48_18;
wire signed[31:0]    reg_activation_48_19;
wire signed[31:0]    reg_activation_48_20;
wire signed[31:0]    reg_activation_48_21;
wire signed[31:0]    reg_activation_48_22;
wire signed[31:0]    reg_activation_48_23;
wire signed[31:0]    reg_activation_48_24;
wire signed[31:0]    reg_activation_48_25;
wire signed[31:0]    reg_activation_48_26;
wire signed[31:0]    reg_activation_48_27;
wire signed[31:0]    reg_activation_48_28;
wire signed[31:0]    reg_activation_48_29;
wire signed[31:0]    reg_activation_48_30;
wire signed[31:0]    reg_activation_48_31;
wire signed[31:0]    reg_activation_48_32;
wire signed[31:0]    reg_activation_48_33;
wire signed[31:0]    reg_activation_48_34;
wire signed[31:0]    reg_activation_48_35;
wire signed[31:0]    reg_activation_48_36;
wire signed[31:0]    reg_activation_48_37;
wire signed[31:0]    reg_activation_48_38;
wire signed[31:0]    reg_activation_48_39;
wire signed[31:0]    reg_activation_48_40;
wire signed[31:0]    reg_activation_48_41;
wire signed[31:0]    reg_activation_48_42;
wire signed[31:0]    reg_activation_48_43;
wire signed[31:0]    reg_activation_48_44;
wire signed[31:0]    reg_activation_48_45;
wire signed[31:0]    reg_activation_48_46;
wire signed[31:0]    reg_activation_48_47;
wire signed[31:0]    reg_activation_48_48;
wire signed[31:0]    reg_activation_48_49;
wire signed[31:0]    reg_activation_48_50;
wire signed[31:0]    reg_activation_48_51;
wire signed[31:0]    reg_activation_48_52;
wire signed[31:0]    reg_activation_48_53;
wire signed[31:0]    reg_activation_48_54;
wire signed[31:0]    reg_activation_48_55;
wire signed[31:0]    reg_activation_48_56;
wire signed[31:0]    reg_activation_48_57;
wire signed[31:0]    reg_activation_48_58;
wire signed[31:0]    reg_activation_48_59;
wire signed[31:0]    reg_activation_48_60;
wire signed[31:0]    reg_activation_48_61;
wire signed[31:0]    reg_activation_48_62;
wire signed[31:0]    reg_activation_48_63;
wire signed[31:0]    reg_activation_49_0;
wire signed[31:0]    reg_activation_49_1;
wire signed[31:0]    reg_activation_49_2;
wire signed[31:0]    reg_activation_49_3;
wire signed[31:0]    reg_activation_49_4;
wire signed[31:0]    reg_activation_49_5;
wire signed[31:0]    reg_activation_49_6;
wire signed[31:0]    reg_activation_49_7;
wire signed[31:0]    reg_activation_49_8;
wire signed[31:0]    reg_activation_49_9;
wire signed[31:0]    reg_activation_49_10;
wire signed[31:0]    reg_activation_49_11;
wire signed[31:0]    reg_activation_49_12;
wire signed[31:0]    reg_activation_49_13;
wire signed[31:0]    reg_activation_49_14;
wire signed[31:0]    reg_activation_49_15;
wire signed[31:0]    reg_activation_49_16;
wire signed[31:0]    reg_activation_49_17;
wire signed[31:0]    reg_activation_49_18;
wire signed[31:0]    reg_activation_49_19;
wire signed[31:0]    reg_activation_49_20;
wire signed[31:0]    reg_activation_49_21;
wire signed[31:0]    reg_activation_49_22;
wire signed[31:0]    reg_activation_49_23;
wire signed[31:0]    reg_activation_49_24;
wire signed[31:0]    reg_activation_49_25;
wire signed[31:0]    reg_activation_49_26;
wire signed[31:0]    reg_activation_49_27;
wire signed[31:0]    reg_activation_49_28;
wire signed[31:0]    reg_activation_49_29;
wire signed[31:0]    reg_activation_49_30;
wire signed[31:0]    reg_activation_49_31;
wire signed[31:0]    reg_activation_49_32;
wire signed[31:0]    reg_activation_49_33;
wire signed[31:0]    reg_activation_49_34;
wire signed[31:0]    reg_activation_49_35;
wire signed[31:0]    reg_activation_49_36;
wire signed[31:0]    reg_activation_49_37;
wire signed[31:0]    reg_activation_49_38;
wire signed[31:0]    reg_activation_49_39;
wire signed[31:0]    reg_activation_49_40;
wire signed[31:0]    reg_activation_49_41;
wire signed[31:0]    reg_activation_49_42;
wire signed[31:0]    reg_activation_49_43;
wire signed[31:0]    reg_activation_49_44;
wire signed[31:0]    reg_activation_49_45;
wire signed[31:0]    reg_activation_49_46;
wire signed[31:0]    reg_activation_49_47;
wire signed[31:0]    reg_activation_49_48;
wire signed[31:0]    reg_activation_49_49;
wire signed[31:0]    reg_activation_49_50;
wire signed[31:0]    reg_activation_49_51;
wire signed[31:0]    reg_activation_49_52;
wire signed[31:0]    reg_activation_49_53;
wire signed[31:0]    reg_activation_49_54;
wire signed[31:0]    reg_activation_49_55;
wire signed[31:0]    reg_activation_49_56;
wire signed[31:0]    reg_activation_49_57;
wire signed[31:0]    reg_activation_49_58;
wire signed[31:0]    reg_activation_49_59;
wire signed[31:0]    reg_activation_49_60;
wire signed[31:0]    reg_activation_49_61;
wire signed[31:0]    reg_activation_49_62;
wire signed[31:0]    reg_activation_49_63;
wire signed[31:0]    reg_activation_50_0;
wire signed[31:0]    reg_activation_50_1;
wire signed[31:0]    reg_activation_50_2;
wire signed[31:0]    reg_activation_50_3;
wire signed[31:0]    reg_activation_50_4;
wire signed[31:0]    reg_activation_50_5;
wire signed[31:0]    reg_activation_50_6;
wire signed[31:0]    reg_activation_50_7;
wire signed[31:0]    reg_activation_50_8;
wire signed[31:0]    reg_activation_50_9;
wire signed[31:0]    reg_activation_50_10;
wire signed[31:0]    reg_activation_50_11;
wire signed[31:0]    reg_activation_50_12;
wire signed[31:0]    reg_activation_50_13;
wire signed[31:0]    reg_activation_50_14;
wire signed[31:0]    reg_activation_50_15;
wire signed[31:0]    reg_activation_50_16;
wire signed[31:0]    reg_activation_50_17;
wire signed[31:0]    reg_activation_50_18;
wire signed[31:0]    reg_activation_50_19;
wire signed[31:0]    reg_activation_50_20;
wire signed[31:0]    reg_activation_50_21;
wire signed[31:0]    reg_activation_50_22;
wire signed[31:0]    reg_activation_50_23;
wire signed[31:0]    reg_activation_50_24;
wire signed[31:0]    reg_activation_50_25;
wire signed[31:0]    reg_activation_50_26;
wire signed[31:0]    reg_activation_50_27;
wire signed[31:0]    reg_activation_50_28;
wire signed[31:0]    reg_activation_50_29;
wire signed[31:0]    reg_activation_50_30;
wire signed[31:0]    reg_activation_50_31;
wire signed[31:0]    reg_activation_50_32;
wire signed[31:0]    reg_activation_50_33;
wire signed[31:0]    reg_activation_50_34;
wire signed[31:0]    reg_activation_50_35;
wire signed[31:0]    reg_activation_50_36;
wire signed[31:0]    reg_activation_50_37;
wire signed[31:0]    reg_activation_50_38;
wire signed[31:0]    reg_activation_50_39;
wire signed[31:0]    reg_activation_50_40;
wire signed[31:0]    reg_activation_50_41;
wire signed[31:0]    reg_activation_50_42;
wire signed[31:0]    reg_activation_50_43;
wire signed[31:0]    reg_activation_50_44;
wire signed[31:0]    reg_activation_50_45;
wire signed[31:0]    reg_activation_50_46;
wire signed[31:0]    reg_activation_50_47;
wire signed[31:0]    reg_activation_50_48;
wire signed[31:0]    reg_activation_50_49;
wire signed[31:0]    reg_activation_50_50;
wire signed[31:0]    reg_activation_50_51;
wire signed[31:0]    reg_activation_50_52;
wire signed[31:0]    reg_activation_50_53;
wire signed[31:0]    reg_activation_50_54;
wire signed[31:0]    reg_activation_50_55;
wire signed[31:0]    reg_activation_50_56;
wire signed[31:0]    reg_activation_50_57;
wire signed[31:0]    reg_activation_50_58;
wire signed[31:0]    reg_activation_50_59;
wire signed[31:0]    reg_activation_50_60;
wire signed[31:0]    reg_activation_50_61;
wire signed[31:0]    reg_activation_50_62;
wire signed[31:0]    reg_activation_50_63;
wire signed[31:0]    reg_activation_51_0;
wire signed[31:0]    reg_activation_51_1;
wire signed[31:0]    reg_activation_51_2;
wire signed[31:0]    reg_activation_51_3;
wire signed[31:0]    reg_activation_51_4;
wire signed[31:0]    reg_activation_51_5;
wire signed[31:0]    reg_activation_51_6;
wire signed[31:0]    reg_activation_51_7;
wire signed[31:0]    reg_activation_51_8;
wire signed[31:0]    reg_activation_51_9;
wire signed[31:0]    reg_activation_51_10;
wire signed[31:0]    reg_activation_51_11;
wire signed[31:0]    reg_activation_51_12;
wire signed[31:0]    reg_activation_51_13;
wire signed[31:0]    reg_activation_51_14;
wire signed[31:0]    reg_activation_51_15;
wire signed[31:0]    reg_activation_51_16;
wire signed[31:0]    reg_activation_51_17;
wire signed[31:0]    reg_activation_51_18;
wire signed[31:0]    reg_activation_51_19;
wire signed[31:0]    reg_activation_51_20;
wire signed[31:0]    reg_activation_51_21;
wire signed[31:0]    reg_activation_51_22;
wire signed[31:0]    reg_activation_51_23;
wire signed[31:0]    reg_activation_51_24;
wire signed[31:0]    reg_activation_51_25;
wire signed[31:0]    reg_activation_51_26;
wire signed[31:0]    reg_activation_51_27;
wire signed[31:0]    reg_activation_51_28;
wire signed[31:0]    reg_activation_51_29;
wire signed[31:0]    reg_activation_51_30;
wire signed[31:0]    reg_activation_51_31;
wire signed[31:0]    reg_activation_51_32;
wire signed[31:0]    reg_activation_51_33;
wire signed[31:0]    reg_activation_51_34;
wire signed[31:0]    reg_activation_51_35;
wire signed[31:0]    reg_activation_51_36;
wire signed[31:0]    reg_activation_51_37;
wire signed[31:0]    reg_activation_51_38;
wire signed[31:0]    reg_activation_51_39;
wire signed[31:0]    reg_activation_51_40;
wire signed[31:0]    reg_activation_51_41;
wire signed[31:0]    reg_activation_51_42;
wire signed[31:0]    reg_activation_51_43;
wire signed[31:0]    reg_activation_51_44;
wire signed[31:0]    reg_activation_51_45;
wire signed[31:0]    reg_activation_51_46;
wire signed[31:0]    reg_activation_51_47;
wire signed[31:0]    reg_activation_51_48;
wire signed[31:0]    reg_activation_51_49;
wire signed[31:0]    reg_activation_51_50;
wire signed[31:0]    reg_activation_51_51;
wire signed[31:0]    reg_activation_51_52;
wire signed[31:0]    reg_activation_51_53;
wire signed[31:0]    reg_activation_51_54;
wire signed[31:0]    reg_activation_51_55;
wire signed[31:0]    reg_activation_51_56;
wire signed[31:0]    reg_activation_51_57;
wire signed[31:0]    reg_activation_51_58;
wire signed[31:0]    reg_activation_51_59;
wire signed[31:0]    reg_activation_51_60;
wire signed[31:0]    reg_activation_51_61;
wire signed[31:0]    reg_activation_51_62;
wire signed[31:0]    reg_activation_51_63;
wire signed[31:0]    reg_activation_52_0;
wire signed[31:0]    reg_activation_52_1;
wire signed[31:0]    reg_activation_52_2;
wire signed[31:0]    reg_activation_52_3;
wire signed[31:0]    reg_activation_52_4;
wire signed[31:0]    reg_activation_52_5;
wire signed[31:0]    reg_activation_52_6;
wire signed[31:0]    reg_activation_52_7;
wire signed[31:0]    reg_activation_52_8;
wire signed[31:0]    reg_activation_52_9;
wire signed[31:0]    reg_activation_52_10;
wire signed[31:0]    reg_activation_52_11;
wire signed[31:0]    reg_activation_52_12;
wire signed[31:0]    reg_activation_52_13;
wire signed[31:0]    reg_activation_52_14;
wire signed[31:0]    reg_activation_52_15;
wire signed[31:0]    reg_activation_52_16;
wire signed[31:0]    reg_activation_52_17;
wire signed[31:0]    reg_activation_52_18;
wire signed[31:0]    reg_activation_52_19;
wire signed[31:0]    reg_activation_52_20;
wire signed[31:0]    reg_activation_52_21;
wire signed[31:0]    reg_activation_52_22;
wire signed[31:0]    reg_activation_52_23;
wire signed[31:0]    reg_activation_52_24;
wire signed[31:0]    reg_activation_52_25;
wire signed[31:0]    reg_activation_52_26;
wire signed[31:0]    reg_activation_52_27;
wire signed[31:0]    reg_activation_52_28;
wire signed[31:0]    reg_activation_52_29;
wire signed[31:0]    reg_activation_52_30;
wire signed[31:0]    reg_activation_52_31;
wire signed[31:0]    reg_activation_52_32;
wire signed[31:0]    reg_activation_52_33;
wire signed[31:0]    reg_activation_52_34;
wire signed[31:0]    reg_activation_52_35;
wire signed[31:0]    reg_activation_52_36;
wire signed[31:0]    reg_activation_52_37;
wire signed[31:0]    reg_activation_52_38;
wire signed[31:0]    reg_activation_52_39;
wire signed[31:0]    reg_activation_52_40;
wire signed[31:0]    reg_activation_52_41;
wire signed[31:0]    reg_activation_52_42;
wire signed[31:0]    reg_activation_52_43;
wire signed[31:0]    reg_activation_52_44;
wire signed[31:0]    reg_activation_52_45;
wire signed[31:0]    reg_activation_52_46;
wire signed[31:0]    reg_activation_52_47;
wire signed[31:0]    reg_activation_52_48;
wire signed[31:0]    reg_activation_52_49;
wire signed[31:0]    reg_activation_52_50;
wire signed[31:0]    reg_activation_52_51;
wire signed[31:0]    reg_activation_52_52;
wire signed[31:0]    reg_activation_52_53;
wire signed[31:0]    reg_activation_52_54;
wire signed[31:0]    reg_activation_52_55;
wire signed[31:0]    reg_activation_52_56;
wire signed[31:0]    reg_activation_52_57;
wire signed[31:0]    reg_activation_52_58;
wire signed[31:0]    reg_activation_52_59;
wire signed[31:0]    reg_activation_52_60;
wire signed[31:0]    reg_activation_52_61;
wire signed[31:0]    reg_activation_52_62;
wire signed[31:0]    reg_activation_52_63;
wire signed[31:0]    reg_activation_53_0;
wire signed[31:0]    reg_activation_53_1;
wire signed[31:0]    reg_activation_53_2;
wire signed[31:0]    reg_activation_53_3;
wire signed[31:0]    reg_activation_53_4;
wire signed[31:0]    reg_activation_53_5;
wire signed[31:0]    reg_activation_53_6;
wire signed[31:0]    reg_activation_53_7;
wire signed[31:0]    reg_activation_53_8;
wire signed[31:0]    reg_activation_53_9;
wire signed[31:0]    reg_activation_53_10;
wire signed[31:0]    reg_activation_53_11;
wire signed[31:0]    reg_activation_53_12;
wire signed[31:0]    reg_activation_53_13;
wire signed[31:0]    reg_activation_53_14;
wire signed[31:0]    reg_activation_53_15;
wire signed[31:0]    reg_activation_53_16;
wire signed[31:0]    reg_activation_53_17;
wire signed[31:0]    reg_activation_53_18;
wire signed[31:0]    reg_activation_53_19;
wire signed[31:0]    reg_activation_53_20;
wire signed[31:0]    reg_activation_53_21;
wire signed[31:0]    reg_activation_53_22;
wire signed[31:0]    reg_activation_53_23;
wire signed[31:0]    reg_activation_53_24;
wire signed[31:0]    reg_activation_53_25;
wire signed[31:0]    reg_activation_53_26;
wire signed[31:0]    reg_activation_53_27;
wire signed[31:0]    reg_activation_53_28;
wire signed[31:0]    reg_activation_53_29;
wire signed[31:0]    reg_activation_53_30;
wire signed[31:0]    reg_activation_53_31;
wire signed[31:0]    reg_activation_53_32;
wire signed[31:0]    reg_activation_53_33;
wire signed[31:0]    reg_activation_53_34;
wire signed[31:0]    reg_activation_53_35;
wire signed[31:0]    reg_activation_53_36;
wire signed[31:0]    reg_activation_53_37;
wire signed[31:0]    reg_activation_53_38;
wire signed[31:0]    reg_activation_53_39;
wire signed[31:0]    reg_activation_53_40;
wire signed[31:0]    reg_activation_53_41;
wire signed[31:0]    reg_activation_53_42;
wire signed[31:0]    reg_activation_53_43;
wire signed[31:0]    reg_activation_53_44;
wire signed[31:0]    reg_activation_53_45;
wire signed[31:0]    reg_activation_53_46;
wire signed[31:0]    reg_activation_53_47;
wire signed[31:0]    reg_activation_53_48;
wire signed[31:0]    reg_activation_53_49;
wire signed[31:0]    reg_activation_53_50;
wire signed[31:0]    reg_activation_53_51;
wire signed[31:0]    reg_activation_53_52;
wire signed[31:0]    reg_activation_53_53;
wire signed[31:0]    reg_activation_53_54;
wire signed[31:0]    reg_activation_53_55;
wire signed[31:0]    reg_activation_53_56;
wire signed[31:0]    reg_activation_53_57;
wire signed[31:0]    reg_activation_53_58;
wire signed[31:0]    reg_activation_53_59;
wire signed[31:0]    reg_activation_53_60;
wire signed[31:0]    reg_activation_53_61;
wire signed[31:0]    reg_activation_53_62;
wire signed[31:0]    reg_activation_53_63;
wire signed[31:0]    reg_activation_54_0;
wire signed[31:0]    reg_activation_54_1;
wire signed[31:0]    reg_activation_54_2;
wire signed[31:0]    reg_activation_54_3;
wire signed[31:0]    reg_activation_54_4;
wire signed[31:0]    reg_activation_54_5;
wire signed[31:0]    reg_activation_54_6;
wire signed[31:0]    reg_activation_54_7;
wire signed[31:0]    reg_activation_54_8;
wire signed[31:0]    reg_activation_54_9;
wire signed[31:0]    reg_activation_54_10;
wire signed[31:0]    reg_activation_54_11;
wire signed[31:0]    reg_activation_54_12;
wire signed[31:0]    reg_activation_54_13;
wire signed[31:0]    reg_activation_54_14;
wire signed[31:0]    reg_activation_54_15;
wire signed[31:0]    reg_activation_54_16;
wire signed[31:0]    reg_activation_54_17;
wire signed[31:0]    reg_activation_54_18;
wire signed[31:0]    reg_activation_54_19;
wire signed[31:0]    reg_activation_54_20;
wire signed[31:0]    reg_activation_54_21;
wire signed[31:0]    reg_activation_54_22;
wire signed[31:0]    reg_activation_54_23;
wire signed[31:0]    reg_activation_54_24;
wire signed[31:0]    reg_activation_54_25;
wire signed[31:0]    reg_activation_54_26;
wire signed[31:0]    reg_activation_54_27;
wire signed[31:0]    reg_activation_54_28;
wire signed[31:0]    reg_activation_54_29;
wire signed[31:0]    reg_activation_54_30;
wire signed[31:0]    reg_activation_54_31;
wire signed[31:0]    reg_activation_54_32;
wire signed[31:0]    reg_activation_54_33;
wire signed[31:0]    reg_activation_54_34;
wire signed[31:0]    reg_activation_54_35;
wire signed[31:0]    reg_activation_54_36;
wire signed[31:0]    reg_activation_54_37;
wire signed[31:0]    reg_activation_54_38;
wire signed[31:0]    reg_activation_54_39;
wire signed[31:0]    reg_activation_54_40;
wire signed[31:0]    reg_activation_54_41;
wire signed[31:0]    reg_activation_54_42;
wire signed[31:0]    reg_activation_54_43;
wire signed[31:0]    reg_activation_54_44;
wire signed[31:0]    reg_activation_54_45;
wire signed[31:0]    reg_activation_54_46;
wire signed[31:0]    reg_activation_54_47;
wire signed[31:0]    reg_activation_54_48;
wire signed[31:0]    reg_activation_54_49;
wire signed[31:0]    reg_activation_54_50;
wire signed[31:0]    reg_activation_54_51;
wire signed[31:0]    reg_activation_54_52;
wire signed[31:0]    reg_activation_54_53;
wire signed[31:0]    reg_activation_54_54;
wire signed[31:0]    reg_activation_54_55;
wire signed[31:0]    reg_activation_54_56;
wire signed[31:0]    reg_activation_54_57;
wire signed[31:0]    reg_activation_54_58;
wire signed[31:0]    reg_activation_54_59;
wire signed[31:0]    reg_activation_54_60;
wire signed[31:0]    reg_activation_54_61;
wire signed[31:0]    reg_activation_54_62;
wire signed[31:0]    reg_activation_54_63;
wire signed[31:0]    reg_activation_55_0;
wire signed[31:0]    reg_activation_55_1;
wire signed[31:0]    reg_activation_55_2;
wire signed[31:0]    reg_activation_55_3;
wire signed[31:0]    reg_activation_55_4;
wire signed[31:0]    reg_activation_55_5;
wire signed[31:0]    reg_activation_55_6;
wire signed[31:0]    reg_activation_55_7;
wire signed[31:0]    reg_activation_55_8;
wire signed[31:0]    reg_activation_55_9;
wire signed[31:0]    reg_activation_55_10;
wire signed[31:0]    reg_activation_55_11;
wire signed[31:0]    reg_activation_55_12;
wire signed[31:0]    reg_activation_55_13;
wire signed[31:0]    reg_activation_55_14;
wire signed[31:0]    reg_activation_55_15;
wire signed[31:0]    reg_activation_55_16;
wire signed[31:0]    reg_activation_55_17;
wire signed[31:0]    reg_activation_55_18;
wire signed[31:0]    reg_activation_55_19;
wire signed[31:0]    reg_activation_55_20;
wire signed[31:0]    reg_activation_55_21;
wire signed[31:0]    reg_activation_55_22;
wire signed[31:0]    reg_activation_55_23;
wire signed[31:0]    reg_activation_55_24;
wire signed[31:0]    reg_activation_55_25;
wire signed[31:0]    reg_activation_55_26;
wire signed[31:0]    reg_activation_55_27;
wire signed[31:0]    reg_activation_55_28;
wire signed[31:0]    reg_activation_55_29;
wire signed[31:0]    reg_activation_55_30;
wire signed[31:0]    reg_activation_55_31;
wire signed[31:0]    reg_activation_55_32;
wire signed[31:0]    reg_activation_55_33;
wire signed[31:0]    reg_activation_55_34;
wire signed[31:0]    reg_activation_55_35;
wire signed[31:0]    reg_activation_55_36;
wire signed[31:0]    reg_activation_55_37;
wire signed[31:0]    reg_activation_55_38;
wire signed[31:0]    reg_activation_55_39;
wire signed[31:0]    reg_activation_55_40;
wire signed[31:0]    reg_activation_55_41;
wire signed[31:0]    reg_activation_55_42;
wire signed[31:0]    reg_activation_55_43;
wire signed[31:0]    reg_activation_55_44;
wire signed[31:0]    reg_activation_55_45;
wire signed[31:0]    reg_activation_55_46;
wire signed[31:0]    reg_activation_55_47;
wire signed[31:0]    reg_activation_55_48;
wire signed[31:0]    reg_activation_55_49;
wire signed[31:0]    reg_activation_55_50;
wire signed[31:0]    reg_activation_55_51;
wire signed[31:0]    reg_activation_55_52;
wire signed[31:0]    reg_activation_55_53;
wire signed[31:0]    reg_activation_55_54;
wire signed[31:0]    reg_activation_55_55;
wire signed[31:0]    reg_activation_55_56;
wire signed[31:0]    reg_activation_55_57;
wire signed[31:0]    reg_activation_55_58;
wire signed[31:0]    reg_activation_55_59;
wire signed[31:0]    reg_activation_55_60;
wire signed[31:0]    reg_activation_55_61;
wire signed[31:0]    reg_activation_55_62;
wire signed[31:0]    reg_activation_55_63;
wire signed[31:0]    reg_activation_56_0;
wire signed[31:0]    reg_activation_56_1;
wire signed[31:0]    reg_activation_56_2;
wire signed[31:0]    reg_activation_56_3;
wire signed[31:0]    reg_activation_56_4;
wire signed[31:0]    reg_activation_56_5;
wire signed[31:0]    reg_activation_56_6;
wire signed[31:0]    reg_activation_56_7;
wire signed[31:0]    reg_activation_56_8;
wire signed[31:0]    reg_activation_56_9;
wire signed[31:0]    reg_activation_56_10;
wire signed[31:0]    reg_activation_56_11;
wire signed[31:0]    reg_activation_56_12;
wire signed[31:0]    reg_activation_56_13;
wire signed[31:0]    reg_activation_56_14;
wire signed[31:0]    reg_activation_56_15;
wire signed[31:0]    reg_activation_56_16;
wire signed[31:0]    reg_activation_56_17;
wire signed[31:0]    reg_activation_56_18;
wire signed[31:0]    reg_activation_56_19;
wire signed[31:0]    reg_activation_56_20;
wire signed[31:0]    reg_activation_56_21;
wire signed[31:0]    reg_activation_56_22;
wire signed[31:0]    reg_activation_56_23;
wire signed[31:0]    reg_activation_56_24;
wire signed[31:0]    reg_activation_56_25;
wire signed[31:0]    reg_activation_56_26;
wire signed[31:0]    reg_activation_56_27;
wire signed[31:0]    reg_activation_56_28;
wire signed[31:0]    reg_activation_56_29;
wire signed[31:0]    reg_activation_56_30;
wire signed[31:0]    reg_activation_56_31;
wire signed[31:0]    reg_activation_56_32;
wire signed[31:0]    reg_activation_56_33;
wire signed[31:0]    reg_activation_56_34;
wire signed[31:0]    reg_activation_56_35;
wire signed[31:0]    reg_activation_56_36;
wire signed[31:0]    reg_activation_56_37;
wire signed[31:0]    reg_activation_56_38;
wire signed[31:0]    reg_activation_56_39;
wire signed[31:0]    reg_activation_56_40;
wire signed[31:0]    reg_activation_56_41;
wire signed[31:0]    reg_activation_56_42;
wire signed[31:0]    reg_activation_56_43;
wire signed[31:0]    reg_activation_56_44;
wire signed[31:0]    reg_activation_56_45;
wire signed[31:0]    reg_activation_56_46;
wire signed[31:0]    reg_activation_56_47;
wire signed[31:0]    reg_activation_56_48;
wire signed[31:0]    reg_activation_56_49;
wire signed[31:0]    reg_activation_56_50;
wire signed[31:0]    reg_activation_56_51;
wire signed[31:0]    reg_activation_56_52;
wire signed[31:0]    reg_activation_56_53;
wire signed[31:0]    reg_activation_56_54;
wire signed[31:0]    reg_activation_56_55;
wire signed[31:0]    reg_activation_56_56;
wire signed[31:0]    reg_activation_56_57;
wire signed[31:0]    reg_activation_56_58;
wire signed[31:0]    reg_activation_56_59;
wire signed[31:0]    reg_activation_56_60;
wire signed[31:0]    reg_activation_56_61;
wire signed[31:0]    reg_activation_56_62;
wire signed[31:0]    reg_activation_56_63;
wire signed[31:0]    reg_activation_57_0;
wire signed[31:0]    reg_activation_57_1;
wire signed[31:0]    reg_activation_57_2;
wire signed[31:0]    reg_activation_57_3;
wire signed[31:0]    reg_activation_57_4;
wire signed[31:0]    reg_activation_57_5;
wire signed[31:0]    reg_activation_57_6;
wire signed[31:0]    reg_activation_57_7;
wire signed[31:0]    reg_activation_57_8;
wire signed[31:0]    reg_activation_57_9;
wire signed[31:0]    reg_activation_57_10;
wire signed[31:0]    reg_activation_57_11;
wire signed[31:0]    reg_activation_57_12;
wire signed[31:0]    reg_activation_57_13;
wire signed[31:0]    reg_activation_57_14;
wire signed[31:0]    reg_activation_57_15;
wire signed[31:0]    reg_activation_57_16;
wire signed[31:0]    reg_activation_57_17;
wire signed[31:0]    reg_activation_57_18;
wire signed[31:0]    reg_activation_57_19;
wire signed[31:0]    reg_activation_57_20;
wire signed[31:0]    reg_activation_57_21;
wire signed[31:0]    reg_activation_57_22;
wire signed[31:0]    reg_activation_57_23;
wire signed[31:0]    reg_activation_57_24;
wire signed[31:0]    reg_activation_57_25;
wire signed[31:0]    reg_activation_57_26;
wire signed[31:0]    reg_activation_57_27;
wire signed[31:0]    reg_activation_57_28;
wire signed[31:0]    reg_activation_57_29;
wire signed[31:0]    reg_activation_57_30;
wire signed[31:0]    reg_activation_57_31;
wire signed[31:0]    reg_activation_57_32;
wire signed[31:0]    reg_activation_57_33;
wire signed[31:0]    reg_activation_57_34;
wire signed[31:0]    reg_activation_57_35;
wire signed[31:0]    reg_activation_57_36;
wire signed[31:0]    reg_activation_57_37;
wire signed[31:0]    reg_activation_57_38;
wire signed[31:0]    reg_activation_57_39;
wire signed[31:0]    reg_activation_57_40;
wire signed[31:0]    reg_activation_57_41;
wire signed[31:0]    reg_activation_57_42;
wire signed[31:0]    reg_activation_57_43;
wire signed[31:0]    reg_activation_57_44;
wire signed[31:0]    reg_activation_57_45;
wire signed[31:0]    reg_activation_57_46;
wire signed[31:0]    reg_activation_57_47;
wire signed[31:0]    reg_activation_57_48;
wire signed[31:0]    reg_activation_57_49;
wire signed[31:0]    reg_activation_57_50;
wire signed[31:0]    reg_activation_57_51;
wire signed[31:0]    reg_activation_57_52;
wire signed[31:0]    reg_activation_57_53;
wire signed[31:0]    reg_activation_57_54;
wire signed[31:0]    reg_activation_57_55;
wire signed[31:0]    reg_activation_57_56;
wire signed[31:0]    reg_activation_57_57;
wire signed[31:0]    reg_activation_57_58;
wire signed[31:0]    reg_activation_57_59;
wire signed[31:0]    reg_activation_57_60;
wire signed[31:0]    reg_activation_57_61;
wire signed[31:0]    reg_activation_57_62;
wire signed[31:0]    reg_activation_57_63;
wire signed[31:0]    reg_activation_58_0;
wire signed[31:0]    reg_activation_58_1;
wire signed[31:0]    reg_activation_58_2;
wire signed[31:0]    reg_activation_58_3;
wire signed[31:0]    reg_activation_58_4;
wire signed[31:0]    reg_activation_58_5;
wire signed[31:0]    reg_activation_58_6;
wire signed[31:0]    reg_activation_58_7;
wire signed[31:0]    reg_activation_58_8;
wire signed[31:0]    reg_activation_58_9;
wire signed[31:0]    reg_activation_58_10;
wire signed[31:0]    reg_activation_58_11;
wire signed[31:0]    reg_activation_58_12;
wire signed[31:0]    reg_activation_58_13;
wire signed[31:0]    reg_activation_58_14;
wire signed[31:0]    reg_activation_58_15;
wire signed[31:0]    reg_activation_58_16;
wire signed[31:0]    reg_activation_58_17;
wire signed[31:0]    reg_activation_58_18;
wire signed[31:0]    reg_activation_58_19;
wire signed[31:0]    reg_activation_58_20;
wire signed[31:0]    reg_activation_58_21;
wire signed[31:0]    reg_activation_58_22;
wire signed[31:0]    reg_activation_58_23;
wire signed[31:0]    reg_activation_58_24;
wire signed[31:0]    reg_activation_58_25;
wire signed[31:0]    reg_activation_58_26;
wire signed[31:0]    reg_activation_58_27;
wire signed[31:0]    reg_activation_58_28;
wire signed[31:0]    reg_activation_58_29;
wire signed[31:0]    reg_activation_58_30;
wire signed[31:0]    reg_activation_58_31;
wire signed[31:0]    reg_activation_58_32;
wire signed[31:0]    reg_activation_58_33;
wire signed[31:0]    reg_activation_58_34;
wire signed[31:0]    reg_activation_58_35;
wire signed[31:0]    reg_activation_58_36;
wire signed[31:0]    reg_activation_58_37;
wire signed[31:0]    reg_activation_58_38;
wire signed[31:0]    reg_activation_58_39;
wire signed[31:0]    reg_activation_58_40;
wire signed[31:0]    reg_activation_58_41;
wire signed[31:0]    reg_activation_58_42;
wire signed[31:0]    reg_activation_58_43;
wire signed[31:0]    reg_activation_58_44;
wire signed[31:0]    reg_activation_58_45;
wire signed[31:0]    reg_activation_58_46;
wire signed[31:0]    reg_activation_58_47;
wire signed[31:0]    reg_activation_58_48;
wire signed[31:0]    reg_activation_58_49;
wire signed[31:0]    reg_activation_58_50;
wire signed[31:0]    reg_activation_58_51;
wire signed[31:0]    reg_activation_58_52;
wire signed[31:0]    reg_activation_58_53;
wire signed[31:0]    reg_activation_58_54;
wire signed[31:0]    reg_activation_58_55;
wire signed[31:0]    reg_activation_58_56;
wire signed[31:0]    reg_activation_58_57;
wire signed[31:0]    reg_activation_58_58;
wire signed[31:0]    reg_activation_58_59;
wire signed[31:0]    reg_activation_58_60;
wire signed[31:0]    reg_activation_58_61;
wire signed[31:0]    reg_activation_58_62;
wire signed[31:0]    reg_activation_58_63;
wire signed[31:0]    reg_activation_59_0;
wire signed[31:0]    reg_activation_59_1;
wire signed[31:0]    reg_activation_59_2;
wire signed[31:0]    reg_activation_59_3;
wire signed[31:0]    reg_activation_59_4;
wire signed[31:0]    reg_activation_59_5;
wire signed[31:0]    reg_activation_59_6;
wire signed[31:0]    reg_activation_59_7;
wire signed[31:0]    reg_activation_59_8;
wire signed[31:0]    reg_activation_59_9;
wire signed[31:0]    reg_activation_59_10;
wire signed[31:0]    reg_activation_59_11;
wire signed[31:0]    reg_activation_59_12;
wire signed[31:0]    reg_activation_59_13;
wire signed[31:0]    reg_activation_59_14;
wire signed[31:0]    reg_activation_59_15;
wire signed[31:0]    reg_activation_59_16;
wire signed[31:0]    reg_activation_59_17;
wire signed[31:0]    reg_activation_59_18;
wire signed[31:0]    reg_activation_59_19;
wire signed[31:0]    reg_activation_59_20;
wire signed[31:0]    reg_activation_59_21;
wire signed[31:0]    reg_activation_59_22;
wire signed[31:0]    reg_activation_59_23;
wire signed[31:0]    reg_activation_59_24;
wire signed[31:0]    reg_activation_59_25;
wire signed[31:0]    reg_activation_59_26;
wire signed[31:0]    reg_activation_59_27;
wire signed[31:0]    reg_activation_59_28;
wire signed[31:0]    reg_activation_59_29;
wire signed[31:0]    reg_activation_59_30;
wire signed[31:0]    reg_activation_59_31;
wire signed[31:0]    reg_activation_59_32;
wire signed[31:0]    reg_activation_59_33;
wire signed[31:0]    reg_activation_59_34;
wire signed[31:0]    reg_activation_59_35;
wire signed[31:0]    reg_activation_59_36;
wire signed[31:0]    reg_activation_59_37;
wire signed[31:0]    reg_activation_59_38;
wire signed[31:0]    reg_activation_59_39;
wire signed[31:0]    reg_activation_59_40;
wire signed[31:0]    reg_activation_59_41;
wire signed[31:0]    reg_activation_59_42;
wire signed[31:0]    reg_activation_59_43;
wire signed[31:0]    reg_activation_59_44;
wire signed[31:0]    reg_activation_59_45;
wire signed[31:0]    reg_activation_59_46;
wire signed[31:0]    reg_activation_59_47;
wire signed[31:0]    reg_activation_59_48;
wire signed[31:0]    reg_activation_59_49;
wire signed[31:0]    reg_activation_59_50;
wire signed[31:0]    reg_activation_59_51;
wire signed[31:0]    reg_activation_59_52;
wire signed[31:0]    reg_activation_59_53;
wire signed[31:0]    reg_activation_59_54;
wire signed[31:0]    reg_activation_59_55;
wire signed[31:0]    reg_activation_59_56;
wire signed[31:0]    reg_activation_59_57;
wire signed[31:0]    reg_activation_59_58;
wire signed[31:0]    reg_activation_59_59;
wire signed[31:0]    reg_activation_59_60;
wire signed[31:0]    reg_activation_59_61;
wire signed[31:0]    reg_activation_59_62;
wire signed[31:0]    reg_activation_59_63;
wire signed[31:0]    reg_activation_60_0;
wire signed[31:0]    reg_activation_60_1;
wire signed[31:0]    reg_activation_60_2;
wire signed[31:0]    reg_activation_60_3;
wire signed[31:0]    reg_activation_60_4;
wire signed[31:0]    reg_activation_60_5;
wire signed[31:0]    reg_activation_60_6;
wire signed[31:0]    reg_activation_60_7;
wire signed[31:0]    reg_activation_60_8;
wire signed[31:0]    reg_activation_60_9;
wire signed[31:0]    reg_activation_60_10;
wire signed[31:0]    reg_activation_60_11;
wire signed[31:0]    reg_activation_60_12;
wire signed[31:0]    reg_activation_60_13;
wire signed[31:0]    reg_activation_60_14;
wire signed[31:0]    reg_activation_60_15;
wire signed[31:0]    reg_activation_60_16;
wire signed[31:0]    reg_activation_60_17;
wire signed[31:0]    reg_activation_60_18;
wire signed[31:0]    reg_activation_60_19;
wire signed[31:0]    reg_activation_60_20;
wire signed[31:0]    reg_activation_60_21;
wire signed[31:0]    reg_activation_60_22;
wire signed[31:0]    reg_activation_60_23;
wire signed[31:0]    reg_activation_60_24;
wire signed[31:0]    reg_activation_60_25;
wire signed[31:0]    reg_activation_60_26;
wire signed[31:0]    reg_activation_60_27;
wire signed[31:0]    reg_activation_60_28;
wire signed[31:0]    reg_activation_60_29;
wire signed[31:0]    reg_activation_60_30;
wire signed[31:0]    reg_activation_60_31;
wire signed[31:0]    reg_activation_60_32;
wire signed[31:0]    reg_activation_60_33;
wire signed[31:0]    reg_activation_60_34;
wire signed[31:0]    reg_activation_60_35;
wire signed[31:0]    reg_activation_60_36;
wire signed[31:0]    reg_activation_60_37;
wire signed[31:0]    reg_activation_60_38;
wire signed[31:0]    reg_activation_60_39;
wire signed[31:0]    reg_activation_60_40;
wire signed[31:0]    reg_activation_60_41;
wire signed[31:0]    reg_activation_60_42;
wire signed[31:0]    reg_activation_60_43;
wire signed[31:0]    reg_activation_60_44;
wire signed[31:0]    reg_activation_60_45;
wire signed[31:0]    reg_activation_60_46;
wire signed[31:0]    reg_activation_60_47;
wire signed[31:0]    reg_activation_60_48;
wire signed[31:0]    reg_activation_60_49;
wire signed[31:0]    reg_activation_60_50;
wire signed[31:0]    reg_activation_60_51;
wire signed[31:0]    reg_activation_60_52;
wire signed[31:0]    reg_activation_60_53;
wire signed[31:0]    reg_activation_60_54;
wire signed[31:0]    reg_activation_60_55;
wire signed[31:0]    reg_activation_60_56;
wire signed[31:0]    reg_activation_60_57;
wire signed[31:0]    reg_activation_60_58;
wire signed[31:0]    reg_activation_60_59;
wire signed[31:0]    reg_activation_60_60;
wire signed[31:0]    reg_activation_60_61;
wire signed[31:0]    reg_activation_60_62;
wire signed[31:0]    reg_activation_60_63;
wire signed[31:0]    reg_activation_61_0;
wire signed[31:0]    reg_activation_61_1;
wire signed[31:0]    reg_activation_61_2;
wire signed[31:0]    reg_activation_61_3;
wire signed[31:0]    reg_activation_61_4;
wire signed[31:0]    reg_activation_61_5;
wire signed[31:0]    reg_activation_61_6;
wire signed[31:0]    reg_activation_61_7;
wire signed[31:0]    reg_activation_61_8;
wire signed[31:0]    reg_activation_61_9;
wire signed[31:0]    reg_activation_61_10;
wire signed[31:0]    reg_activation_61_11;
wire signed[31:0]    reg_activation_61_12;
wire signed[31:0]    reg_activation_61_13;
wire signed[31:0]    reg_activation_61_14;
wire signed[31:0]    reg_activation_61_15;
wire signed[31:0]    reg_activation_61_16;
wire signed[31:0]    reg_activation_61_17;
wire signed[31:0]    reg_activation_61_18;
wire signed[31:0]    reg_activation_61_19;
wire signed[31:0]    reg_activation_61_20;
wire signed[31:0]    reg_activation_61_21;
wire signed[31:0]    reg_activation_61_22;
wire signed[31:0]    reg_activation_61_23;
wire signed[31:0]    reg_activation_61_24;
wire signed[31:0]    reg_activation_61_25;
wire signed[31:0]    reg_activation_61_26;
wire signed[31:0]    reg_activation_61_27;
wire signed[31:0]    reg_activation_61_28;
wire signed[31:0]    reg_activation_61_29;
wire signed[31:0]    reg_activation_61_30;
wire signed[31:0]    reg_activation_61_31;
wire signed[31:0]    reg_activation_61_32;
wire signed[31:0]    reg_activation_61_33;
wire signed[31:0]    reg_activation_61_34;
wire signed[31:0]    reg_activation_61_35;
wire signed[31:0]    reg_activation_61_36;
wire signed[31:0]    reg_activation_61_37;
wire signed[31:0]    reg_activation_61_38;
wire signed[31:0]    reg_activation_61_39;
wire signed[31:0]    reg_activation_61_40;
wire signed[31:0]    reg_activation_61_41;
wire signed[31:0]    reg_activation_61_42;
wire signed[31:0]    reg_activation_61_43;
wire signed[31:0]    reg_activation_61_44;
wire signed[31:0]    reg_activation_61_45;
wire signed[31:0]    reg_activation_61_46;
wire signed[31:0]    reg_activation_61_47;
wire signed[31:0]    reg_activation_61_48;
wire signed[31:0]    reg_activation_61_49;
wire signed[31:0]    reg_activation_61_50;
wire signed[31:0]    reg_activation_61_51;
wire signed[31:0]    reg_activation_61_52;
wire signed[31:0]    reg_activation_61_53;
wire signed[31:0]    reg_activation_61_54;
wire signed[31:0]    reg_activation_61_55;
wire signed[31:0]    reg_activation_61_56;
wire signed[31:0]    reg_activation_61_57;
wire signed[31:0]    reg_activation_61_58;
wire signed[31:0]    reg_activation_61_59;
wire signed[31:0]    reg_activation_61_60;
wire signed[31:0]    reg_activation_61_61;
wire signed[31:0]    reg_activation_61_62;
wire signed[31:0]    reg_activation_61_63;
wire signed[31:0]    reg_activation_62_0;
wire signed[31:0]    reg_activation_62_1;
wire signed[31:0]    reg_activation_62_2;
wire signed[31:0]    reg_activation_62_3;
wire signed[31:0]    reg_activation_62_4;
wire signed[31:0]    reg_activation_62_5;
wire signed[31:0]    reg_activation_62_6;
wire signed[31:0]    reg_activation_62_7;
wire signed[31:0]    reg_activation_62_8;
wire signed[31:0]    reg_activation_62_9;
wire signed[31:0]    reg_activation_62_10;
wire signed[31:0]    reg_activation_62_11;
wire signed[31:0]    reg_activation_62_12;
wire signed[31:0]    reg_activation_62_13;
wire signed[31:0]    reg_activation_62_14;
wire signed[31:0]    reg_activation_62_15;
wire signed[31:0]    reg_activation_62_16;
wire signed[31:0]    reg_activation_62_17;
wire signed[31:0]    reg_activation_62_18;
wire signed[31:0]    reg_activation_62_19;
wire signed[31:0]    reg_activation_62_20;
wire signed[31:0]    reg_activation_62_21;
wire signed[31:0]    reg_activation_62_22;
wire signed[31:0]    reg_activation_62_23;
wire signed[31:0]    reg_activation_62_24;
wire signed[31:0]    reg_activation_62_25;
wire signed[31:0]    reg_activation_62_26;
wire signed[31:0]    reg_activation_62_27;
wire signed[31:0]    reg_activation_62_28;
wire signed[31:0]    reg_activation_62_29;
wire signed[31:0]    reg_activation_62_30;
wire signed[31:0]    reg_activation_62_31;
wire signed[31:0]    reg_activation_62_32;
wire signed[31:0]    reg_activation_62_33;
wire signed[31:0]    reg_activation_62_34;
wire signed[31:0]    reg_activation_62_35;
wire signed[31:0]    reg_activation_62_36;
wire signed[31:0]    reg_activation_62_37;
wire signed[31:0]    reg_activation_62_38;
wire signed[31:0]    reg_activation_62_39;
wire signed[31:0]    reg_activation_62_40;
wire signed[31:0]    reg_activation_62_41;
wire signed[31:0]    reg_activation_62_42;
wire signed[31:0]    reg_activation_62_43;
wire signed[31:0]    reg_activation_62_44;
wire signed[31:0]    reg_activation_62_45;
wire signed[31:0]    reg_activation_62_46;
wire signed[31:0]    reg_activation_62_47;
wire signed[31:0]    reg_activation_62_48;
wire signed[31:0]    reg_activation_62_49;
wire signed[31:0]    reg_activation_62_50;
wire signed[31:0]    reg_activation_62_51;
wire signed[31:0]    reg_activation_62_52;
wire signed[31:0]    reg_activation_62_53;
wire signed[31:0]    reg_activation_62_54;
wire signed[31:0]    reg_activation_62_55;
wire signed[31:0]    reg_activation_62_56;
wire signed[31:0]    reg_activation_62_57;
wire signed[31:0]    reg_activation_62_58;
wire signed[31:0]    reg_activation_62_59;
wire signed[31:0]    reg_activation_62_60;
wire signed[31:0]    reg_activation_62_61;
wire signed[31:0]    reg_activation_62_62;
wire signed[31:0]    reg_activation_62_63;
wire signed[31:0]    reg_activation_63_0;
wire signed[31:0]    reg_activation_63_1;
wire signed[31:0]    reg_activation_63_2;
wire signed[31:0]    reg_activation_63_3;
wire signed[31:0]    reg_activation_63_4;
wire signed[31:0]    reg_activation_63_5;
wire signed[31:0]    reg_activation_63_6;
wire signed[31:0]    reg_activation_63_7;
wire signed[31:0]    reg_activation_63_8;
wire signed[31:0]    reg_activation_63_9;
wire signed[31:0]    reg_activation_63_10;
wire signed[31:0]    reg_activation_63_11;
wire signed[31:0]    reg_activation_63_12;
wire signed[31:0]    reg_activation_63_13;
wire signed[31:0]    reg_activation_63_14;
wire signed[31:0]    reg_activation_63_15;
wire signed[31:0]    reg_activation_63_16;
wire signed[31:0]    reg_activation_63_17;
wire signed[31:0]    reg_activation_63_18;
wire signed[31:0]    reg_activation_63_19;
wire signed[31:0]    reg_activation_63_20;
wire signed[31:0]    reg_activation_63_21;
wire signed[31:0]    reg_activation_63_22;
wire signed[31:0]    reg_activation_63_23;
wire signed[31:0]    reg_activation_63_24;
wire signed[31:0]    reg_activation_63_25;
wire signed[31:0]    reg_activation_63_26;
wire signed[31:0]    reg_activation_63_27;
wire signed[31:0]    reg_activation_63_28;
wire signed[31:0]    reg_activation_63_29;
wire signed[31:0]    reg_activation_63_30;
wire signed[31:0]    reg_activation_63_31;
wire signed[31:0]    reg_activation_63_32;
wire signed[31:0]    reg_activation_63_33;
wire signed[31:0]    reg_activation_63_34;
wire signed[31:0]    reg_activation_63_35;
wire signed[31:0]    reg_activation_63_36;
wire signed[31:0]    reg_activation_63_37;
wire signed[31:0]    reg_activation_63_38;
wire signed[31:0]    reg_activation_63_39;
wire signed[31:0]    reg_activation_63_40;
wire signed[31:0]    reg_activation_63_41;
wire signed[31:0]    reg_activation_63_42;
wire signed[31:0]    reg_activation_63_43;
wire signed[31:0]    reg_activation_63_44;
wire signed[31:0]    reg_activation_63_45;
wire signed[31:0]    reg_activation_63_46;
wire signed[31:0]    reg_activation_63_47;
wire signed[31:0]    reg_activation_63_48;
wire signed[31:0]    reg_activation_63_49;
wire signed[31:0]    reg_activation_63_50;
wire signed[31:0]    reg_activation_63_51;
wire signed[31:0]    reg_activation_63_52;
wire signed[31:0]    reg_activation_63_53;
wire signed[31:0]    reg_activation_63_54;
wire signed[31:0]    reg_activation_63_55;
wire signed[31:0]    reg_activation_63_56;
wire signed[31:0]    reg_activation_63_57;
wire signed[31:0]    reg_activation_63_58;
wire signed[31:0]    reg_activation_63_59;
wire signed[31:0]    reg_activation_63_60;
wire signed[31:0]    reg_activation_63_61;
wire signed[31:0]    reg_activation_63_62;
wire signed[31:0]    reg_activation_63_63;
wire signed[31:0]    reg_weight_0_0;
wire signed[31:0]    reg_psum_0_0;
wire signed[31:0]    reg_weight_0_1;
wire signed[31:0]    reg_psum_0_1;
wire signed[31:0]    reg_weight_0_2;
wire signed[31:0]    reg_psum_0_2;
wire signed[31:0]    reg_weight_0_3;
wire signed[31:0]    reg_psum_0_3;
wire signed[31:0]    reg_weight_0_4;
wire signed[31:0]    reg_psum_0_4;
wire signed[31:0]    reg_weight_0_5;
wire signed[31:0]    reg_psum_0_5;
wire signed[31:0]    reg_weight_0_6;
wire signed[31:0]    reg_psum_0_6;
wire signed[31:0]    reg_weight_0_7;
wire signed[31:0]    reg_psum_0_7;
wire signed[31:0]    reg_weight_0_8;
wire signed[31:0]    reg_psum_0_8;
wire signed[31:0]    reg_weight_0_9;
wire signed[31:0]    reg_psum_0_9;
wire signed[31:0]    reg_weight_0_10;
wire signed[31:0]    reg_psum_0_10;
wire signed[31:0]    reg_weight_0_11;
wire signed[31:0]    reg_psum_0_11;
wire signed[31:0]    reg_weight_0_12;
wire signed[31:0]    reg_psum_0_12;
wire signed[31:0]    reg_weight_0_13;
wire signed[31:0]    reg_psum_0_13;
wire signed[31:0]    reg_weight_0_14;
wire signed[31:0]    reg_psum_0_14;
wire signed[31:0]    reg_weight_0_15;
wire signed[31:0]    reg_psum_0_15;
wire signed[31:0]    reg_weight_0_16;
wire signed[31:0]    reg_psum_0_16;
wire signed[31:0]    reg_weight_0_17;
wire signed[31:0]    reg_psum_0_17;
wire signed[31:0]    reg_weight_0_18;
wire signed[31:0]    reg_psum_0_18;
wire signed[31:0]    reg_weight_0_19;
wire signed[31:0]    reg_psum_0_19;
wire signed[31:0]    reg_weight_0_20;
wire signed[31:0]    reg_psum_0_20;
wire signed[31:0]    reg_weight_0_21;
wire signed[31:0]    reg_psum_0_21;
wire signed[31:0]    reg_weight_0_22;
wire signed[31:0]    reg_psum_0_22;
wire signed[31:0]    reg_weight_0_23;
wire signed[31:0]    reg_psum_0_23;
wire signed[31:0]    reg_weight_0_24;
wire signed[31:0]    reg_psum_0_24;
wire signed[31:0]    reg_weight_0_25;
wire signed[31:0]    reg_psum_0_25;
wire signed[31:0]    reg_weight_0_26;
wire signed[31:0]    reg_psum_0_26;
wire signed[31:0]    reg_weight_0_27;
wire signed[31:0]    reg_psum_0_27;
wire signed[31:0]    reg_weight_0_28;
wire signed[31:0]    reg_psum_0_28;
wire signed[31:0]    reg_weight_0_29;
wire signed[31:0]    reg_psum_0_29;
wire signed[31:0]    reg_weight_0_30;
wire signed[31:0]    reg_psum_0_30;
wire signed[31:0]    reg_weight_0_31;
wire signed[31:0]    reg_psum_0_31;
wire signed[31:0]    reg_weight_0_32;
wire signed[31:0]    reg_psum_0_32;
wire signed[31:0]    reg_weight_0_33;
wire signed[31:0]    reg_psum_0_33;
wire signed[31:0]    reg_weight_0_34;
wire signed[31:0]    reg_psum_0_34;
wire signed[31:0]    reg_weight_0_35;
wire signed[31:0]    reg_psum_0_35;
wire signed[31:0]    reg_weight_0_36;
wire signed[31:0]    reg_psum_0_36;
wire signed[31:0]    reg_weight_0_37;
wire signed[31:0]    reg_psum_0_37;
wire signed[31:0]    reg_weight_0_38;
wire signed[31:0]    reg_psum_0_38;
wire signed[31:0]    reg_weight_0_39;
wire signed[31:0]    reg_psum_0_39;
wire signed[31:0]    reg_weight_0_40;
wire signed[31:0]    reg_psum_0_40;
wire signed[31:0]    reg_weight_0_41;
wire signed[31:0]    reg_psum_0_41;
wire signed[31:0]    reg_weight_0_42;
wire signed[31:0]    reg_psum_0_42;
wire signed[31:0]    reg_weight_0_43;
wire signed[31:0]    reg_psum_0_43;
wire signed[31:0]    reg_weight_0_44;
wire signed[31:0]    reg_psum_0_44;
wire signed[31:0]    reg_weight_0_45;
wire signed[31:0]    reg_psum_0_45;
wire signed[31:0]    reg_weight_0_46;
wire signed[31:0]    reg_psum_0_46;
wire signed[31:0]    reg_weight_0_47;
wire signed[31:0]    reg_psum_0_47;
wire signed[31:0]    reg_weight_0_48;
wire signed[31:0]    reg_psum_0_48;
wire signed[31:0]    reg_weight_0_49;
wire signed[31:0]    reg_psum_0_49;
wire signed[31:0]    reg_weight_0_50;
wire signed[31:0]    reg_psum_0_50;
wire signed[31:0]    reg_weight_0_51;
wire signed[31:0]    reg_psum_0_51;
wire signed[31:0]    reg_weight_0_52;
wire signed[31:0]    reg_psum_0_52;
wire signed[31:0]    reg_weight_0_53;
wire signed[31:0]    reg_psum_0_53;
wire signed[31:0]    reg_weight_0_54;
wire signed[31:0]    reg_psum_0_54;
wire signed[31:0]    reg_weight_0_55;
wire signed[31:0]    reg_psum_0_55;
wire signed[31:0]    reg_weight_0_56;
wire signed[31:0]    reg_psum_0_56;
wire signed[31:0]    reg_weight_0_57;
wire signed[31:0]    reg_psum_0_57;
wire signed[31:0]    reg_weight_0_58;
wire signed[31:0]    reg_psum_0_58;
wire signed[31:0]    reg_weight_0_59;
wire signed[31:0]    reg_psum_0_59;
wire signed[31:0]    reg_weight_0_60;
wire signed[31:0]    reg_psum_0_60;
wire signed[31:0]    reg_weight_0_61;
wire signed[31:0]    reg_psum_0_61;
wire signed[31:0]    reg_weight_0_62;
wire signed[31:0]    reg_psum_0_62;
wire signed[31:0]    reg_weight_0_63;
wire signed[31:0]    reg_psum_0_63;
wire signed[31:0]    reg_weight_1_0;
wire signed[31:0]    reg_psum_1_0;
wire signed[31:0]    reg_weight_1_1;
wire signed[31:0]    reg_psum_1_1;
wire signed[31:0]    reg_weight_1_2;
wire signed[31:0]    reg_psum_1_2;
wire signed[31:0]    reg_weight_1_3;
wire signed[31:0]    reg_psum_1_3;
wire signed[31:0]    reg_weight_1_4;
wire signed[31:0]    reg_psum_1_4;
wire signed[31:0]    reg_weight_1_5;
wire signed[31:0]    reg_psum_1_5;
wire signed[31:0]    reg_weight_1_6;
wire signed[31:0]    reg_psum_1_6;
wire signed[31:0]    reg_weight_1_7;
wire signed[31:0]    reg_psum_1_7;
wire signed[31:0]    reg_weight_1_8;
wire signed[31:0]    reg_psum_1_8;
wire signed[31:0]    reg_weight_1_9;
wire signed[31:0]    reg_psum_1_9;
wire signed[31:0]    reg_weight_1_10;
wire signed[31:0]    reg_psum_1_10;
wire signed[31:0]    reg_weight_1_11;
wire signed[31:0]    reg_psum_1_11;
wire signed[31:0]    reg_weight_1_12;
wire signed[31:0]    reg_psum_1_12;
wire signed[31:0]    reg_weight_1_13;
wire signed[31:0]    reg_psum_1_13;
wire signed[31:0]    reg_weight_1_14;
wire signed[31:0]    reg_psum_1_14;
wire signed[31:0]    reg_weight_1_15;
wire signed[31:0]    reg_psum_1_15;
wire signed[31:0]    reg_weight_1_16;
wire signed[31:0]    reg_psum_1_16;
wire signed[31:0]    reg_weight_1_17;
wire signed[31:0]    reg_psum_1_17;
wire signed[31:0]    reg_weight_1_18;
wire signed[31:0]    reg_psum_1_18;
wire signed[31:0]    reg_weight_1_19;
wire signed[31:0]    reg_psum_1_19;
wire signed[31:0]    reg_weight_1_20;
wire signed[31:0]    reg_psum_1_20;
wire signed[31:0]    reg_weight_1_21;
wire signed[31:0]    reg_psum_1_21;
wire signed[31:0]    reg_weight_1_22;
wire signed[31:0]    reg_psum_1_22;
wire signed[31:0]    reg_weight_1_23;
wire signed[31:0]    reg_psum_1_23;
wire signed[31:0]    reg_weight_1_24;
wire signed[31:0]    reg_psum_1_24;
wire signed[31:0]    reg_weight_1_25;
wire signed[31:0]    reg_psum_1_25;
wire signed[31:0]    reg_weight_1_26;
wire signed[31:0]    reg_psum_1_26;
wire signed[31:0]    reg_weight_1_27;
wire signed[31:0]    reg_psum_1_27;
wire signed[31:0]    reg_weight_1_28;
wire signed[31:0]    reg_psum_1_28;
wire signed[31:0]    reg_weight_1_29;
wire signed[31:0]    reg_psum_1_29;
wire signed[31:0]    reg_weight_1_30;
wire signed[31:0]    reg_psum_1_30;
wire signed[31:0]    reg_weight_1_31;
wire signed[31:0]    reg_psum_1_31;
wire signed[31:0]    reg_weight_1_32;
wire signed[31:0]    reg_psum_1_32;
wire signed[31:0]    reg_weight_1_33;
wire signed[31:0]    reg_psum_1_33;
wire signed[31:0]    reg_weight_1_34;
wire signed[31:0]    reg_psum_1_34;
wire signed[31:0]    reg_weight_1_35;
wire signed[31:0]    reg_psum_1_35;
wire signed[31:0]    reg_weight_1_36;
wire signed[31:0]    reg_psum_1_36;
wire signed[31:0]    reg_weight_1_37;
wire signed[31:0]    reg_psum_1_37;
wire signed[31:0]    reg_weight_1_38;
wire signed[31:0]    reg_psum_1_38;
wire signed[31:0]    reg_weight_1_39;
wire signed[31:0]    reg_psum_1_39;
wire signed[31:0]    reg_weight_1_40;
wire signed[31:0]    reg_psum_1_40;
wire signed[31:0]    reg_weight_1_41;
wire signed[31:0]    reg_psum_1_41;
wire signed[31:0]    reg_weight_1_42;
wire signed[31:0]    reg_psum_1_42;
wire signed[31:0]    reg_weight_1_43;
wire signed[31:0]    reg_psum_1_43;
wire signed[31:0]    reg_weight_1_44;
wire signed[31:0]    reg_psum_1_44;
wire signed[31:0]    reg_weight_1_45;
wire signed[31:0]    reg_psum_1_45;
wire signed[31:0]    reg_weight_1_46;
wire signed[31:0]    reg_psum_1_46;
wire signed[31:0]    reg_weight_1_47;
wire signed[31:0]    reg_psum_1_47;
wire signed[31:0]    reg_weight_1_48;
wire signed[31:0]    reg_psum_1_48;
wire signed[31:0]    reg_weight_1_49;
wire signed[31:0]    reg_psum_1_49;
wire signed[31:0]    reg_weight_1_50;
wire signed[31:0]    reg_psum_1_50;
wire signed[31:0]    reg_weight_1_51;
wire signed[31:0]    reg_psum_1_51;
wire signed[31:0]    reg_weight_1_52;
wire signed[31:0]    reg_psum_1_52;
wire signed[31:0]    reg_weight_1_53;
wire signed[31:0]    reg_psum_1_53;
wire signed[31:0]    reg_weight_1_54;
wire signed[31:0]    reg_psum_1_54;
wire signed[31:0]    reg_weight_1_55;
wire signed[31:0]    reg_psum_1_55;
wire signed[31:0]    reg_weight_1_56;
wire signed[31:0]    reg_psum_1_56;
wire signed[31:0]    reg_weight_1_57;
wire signed[31:0]    reg_psum_1_57;
wire signed[31:0]    reg_weight_1_58;
wire signed[31:0]    reg_psum_1_58;
wire signed[31:0]    reg_weight_1_59;
wire signed[31:0]    reg_psum_1_59;
wire signed[31:0]    reg_weight_1_60;
wire signed[31:0]    reg_psum_1_60;
wire signed[31:0]    reg_weight_1_61;
wire signed[31:0]    reg_psum_1_61;
wire signed[31:0]    reg_weight_1_62;
wire signed[31:0]    reg_psum_1_62;
wire signed[31:0]    reg_weight_1_63;
wire signed[31:0]    reg_psum_1_63;
wire signed[31:0]    reg_weight_2_0;
wire signed[31:0]    reg_psum_2_0;
wire signed[31:0]    reg_weight_2_1;
wire signed[31:0]    reg_psum_2_1;
wire signed[31:0]    reg_weight_2_2;
wire signed[31:0]    reg_psum_2_2;
wire signed[31:0]    reg_weight_2_3;
wire signed[31:0]    reg_psum_2_3;
wire signed[31:0]    reg_weight_2_4;
wire signed[31:0]    reg_psum_2_4;
wire signed[31:0]    reg_weight_2_5;
wire signed[31:0]    reg_psum_2_5;
wire signed[31:0]    reg_weight_2_6;
wire signed[31:0]    reg_psum_2_6;
wire signed[31:0]    reg_weight_2_7;
wire signed[31:0]    reg_psum_2_7;
wire signed[31:0]    reg_weight_2_8;
wire signed[31:0]    reg_psum_2_8;
wire signed[31:0]    reg_weight_2_9;
wire signed[31:0]    reg_psum_2_9;
wire signed[31:0]    reg_weight_2_10;
wire signed[31:0]    reg_psum_2_10;
wire signed[31:0]    reg_weight_2_11;
wire signed[31:0]    reg_psum_2_11;
wire signed[31:0]    reg_weight_2_12;
wire signed[31:0]    reg_psum_2_12;
wire signed[31:0]    reg_weight_2_13;
wire signed[31:0]    reg_psum_2_13;
wire signed[31:0]    reg_weight_2_14;
wire signed[31:0]    reg_psum_2_14;
wire signed[31:0]    reg_weight_2_15;
wire signed[31:0]    reg_psum_2_15;
wire signed[31:0]    reg_weight_2_16;
wire signed[31:0]    reg_psum_2_16;
wire signed[31:0]    reg_weight_2_17;
wire signed[31:0]    reg_psum_2_17;
wire signed[31:0]    reg_weight_2_18;
wire signed[31:0]    reg_psum_2_18;
wire signed[31:0]    reg_weight_2_19;
wire signed[31:0]    reg_psum_2_19;
wire signed[31:0]    reg_weight_2_20;
wire signed[31:0]    reg_psum_2_20;
wire signed[31:0]    reg_weight_2_21;
wire signed[31:0]    reg_psum_2_21;
wire signed[31:0]    reg_weight_2_22;
wire signed[31:0]    reg_psum_2_22;
wire signed[31:0]    reg_weight_2_23;
wire signed[31:0]    reg_psum_2_23;
wire signed[31:0]    reg_weight_2_24;
wire signed[31:0]    reg_psum_2_24;
wire signed[31:0]    reg_weight_2_25;
wire signed[31:0]    reg_psum_2_25;
wire signed[31:0]    reg_weight_2_26;
wire signed[31:0]    reg_psum_2_26;
wire signed[31:0]    reg_weight_2_27;
wire signed[31:0]    reg_psum_2_27;
wire signed[31:0]    reg_weight_2_28;
wire signed[31:0]    reg_psum_2_28;
wire signed[31:0]    reg_weight_2_29;
wire signed[31:0]    reg_psum_2_29;
wire signed[31:0]    reg_weight_2_30;
wire signed[31:0]    reg_psum_2_30;
wire signed[31:0]    reg_weight_2_31;
wire signed[31:0]    reg_psum_2_31;
wire signed[31:0]    reg_weight_2_32;
wire signed[31:0]    reg_psum_2_32;
wire signed[31:0]    reg_weight_2_33;
wire signed[31:0]    reg_psum_2_33;
wire signed[31:0]    reg_weight_2_34;
wire signed[31:0]    reg_psum_2_34;
wire signed[31:0]    reg_weight_2_35;
wire signed[31:0]    reg_psum_2_35;
wire signed[31:0]    reg_weight_2_36;
wire signed[31:0]    reg_psum_2_36;
wire signed[31:0]    reg_weight_2_37;
wire signed[31:0]    reg_psum_2_37;
wire signed[31:0]    reg_weight_2_38;
wire signed[31:0]    reg_psum_2_38;
wire signed[31:0]    reg_weight_2_39;
wire signed[31:0]    reg_psum_2_39;
wire signed[31:0]    reg_weight_2_40;
wire signed[31:0]    reg_psum_2_40;
wire signed[31:0]    reg_weight_2_41;
wire signed[31:0]    reg_psum_2_41;
wire signed[31:0]    reg_weight_2_42;
wire signed[31:0]    reg_psum_2_42;
wire signed[31:0]    reg_weight_2_43;
wire signed[31:0]    reg_psum_2_43;
wire signed[31:0]    reg_weight_2_44;
wire signed[31:0]    reg_psum_2_44;
wire signed[31:0]    reg_weight_2_45;
wire signed[31:0]    reg_psum_2_45;
wire signed[31:0]    reg_weight_2_46;
wire signed[31:0]    reg_psum_2_46;
wire signed[31:0]    reg_weight_2_47;
wire signed[31:0]    reg_psum_2_47;
wire signed[31:0]    reg_weight_2_48;
wire signed[31:0]    reg_psum_2_48;
wire signed[31:0]    reg_weight_2_49;
wire signed[31:0]    reg_psum_2_49;
wire signed[31:0]    reg_weight_2_50;
wire signed[31:0]    reg_psum_2_50;
wire signed[31:0]    reg_weight_2_51;
wire signed[31:0]    reg_psum_2_51;
wire signed[31:0]    reg_weight_2_52;
wire signed[31:0]    reg_psum_2_52;
wire signed[31:0]    reg_weight_2_53;
wire signed[31:0]    reg_psum_2_53;
wire signed[31:0]    reg_weight_2_54;
wire signed[31:0]    reg_psum_2_54;
wire signed[31:0]    reg_weight_2_55;
wire signed[31:0]    reg_psum_2_55;
wire signed[31:0]    reg_weight_2_56;
wire signed[31:0]    reg_psum_2_56;
wire signed[31:0]    reg_weight_2_57;
wire signed[31:0]    reg_psum_2_57;
wire signed[31:0]    reg_weight_2_58;
wire signed[31:0]    reg_psum_2_58;
wire signed[31:0]    reg_weight_2_59;
wire signed[31:0]    reg_psum_2_59;
wire signed[31:0]    reg_weight_2_60;
wire signed[31:0]    reg_psum_2_60;
wire signed[31:0]    reg_weight_2_61;
wire signed[31:0]    reg_psum_2_61;
wire signed[31:0]    reg_weight_2_62;
wire signed[31:0]    reg_psum_2_62;
wire signed[31:0]    reg_weight_2_63;
wire signed[31:0]    reg_psum_2_63;
wire signed[31:0]    reg_weight_3_0;
wire signed[31:0]    reg_psum_3_0;
wire signed[31:0]    reg_weight_3_1;
wire signed[31:0]    reg_psum_3_1;
wire signed[31:0]    reg_weight_3_2;
wire signed[31:0]    reg_psum_3_2;
wire signed[31:0]    reg_weight_3_3;
wire signed[31:0]    reg_psum_3_3;
wire signed[31:0]    reg_weight_3_4;
wire signed[31:0]    reg_psum_3_4;
wire signed[31:0]    reg_weight_3_5;
wire signed[31:0]    reg_psum_3_5;
wire signed[31:0]    reg_weight_3_6;
wire signed[31:0]    reg_psum_3_6;
wire signed[31:0]    reg_weight_3_7;
wire signed[31:0]    reg_psum_3_7;
wire signed[31:0]    reg_weight_3_8;
wire signed[31:0]    reg_psum_3_8;
wire signed[31:0]    reg_weight_3_9;
wire signed[31:0]    reg_psum_3_9;
wire signed[31:0]    reg_weight_3_10;
wire signed[31:0]    reg_psum_3_10;
wire signed[31:0]    reg_weight_3_11;
wire signed[31:0]    reg_psum_3_11;
wire signed[31:0]    reg_weight_3_12;
wire signed[31:0]    reg_psum_3_12;
wire signed[31:0]    reg_weight_3_13;
wire signed[31:0]    reg_psum_3_13;
wire signed[31:0]    reg_weight_3_14;
wire signed[31:0]    reg_psum_3_14;
wire signed[31:0]    reg_weight_3_15;
wire signed[31:0]    reg_psum_3_15;
wire signed[31:0]    reg_weight_3_16;
wire signed[31:0]    reg_psum_3_16;
wire signed[31:0]    reg_weight_3_17;
wire signed[31:0]    reg_psum_3_17;
wire signed[31:0]    reg_weight_3_18;
wire signed[31:0]    reg_psum_3_18;
wire signed[31:0]    reg_weight_3_19;
wire signed[31:0]    reg_psum_3_19;
wire signed[31:0]    reg_weight_3_20;
wire signed[31:0]    reg_psum_3_20;
wire signed[31:0]    reg_weight_3_21;
wire signed[31:0]    reg_psum_3_21;
wire signed[31:0]    reg_weight_3_22;
wire signed[31:0]    reg_psum_3_22;
wire signed[31:0]    reg_weight_3_23;
wire signed[31:0]    reg_psum_3_23;
wire signed[31:0]    reg_weight_3_24;
wire signed[31:0]    reg_psum_3_24;
wire signed[31:0]    reg_weight_3_25;
wire signed[31:0]    reg_psum_3_25;
wire signed[31:0]    reg_weight_3_26;
wire signed[31:0]    reg_psum_3_26;
wire signed[31:0]    reg_weight_3_27;
wire signed[31:0]    reg_psum_3_27;
wire signed[31:0]    reg_weight_3_28;
wire signed[31:0]    reg_psum_3_28;
wire signed[31:0]    reg_weight_3_29;
wire signed[31:0]    reg_psum_3_29;
wire signed[31:0]    reg_weight_3_30;
wire signed[31:0]    reg_psum_3_30;
wire signed[31:0]    reg_weight_3_31;
wire signed[31:0]    reg_psum_3_31;
wire signed[31:0]    reg_weight_3_32;
wire signed[31:0]    reg_psum_3_32;
wire signed[31:0]    reg_weight_3_33;
wire signed[31:0]    reg_psum_3_33;
wire signed[31:0]    reg_weight_3_34;
wire signed[31:0]    reg_psum_3_34;
wire signed[31:0]    reg_weight_3_35;
wire signed[31:0]    reg_psum_3_35;
wire signed[31:0]    reg_weight_3_36;
wire signed[31:0]    reg_psum_3_36;
wire signed[31:0]    reg_weight_3_37;
wire signed[31:0]    reg_psum_3_37;
wire signed[31:0]    reg_weight_3_38;
wire signed[31:0]    reg_psum_3_38;
wire signed[31:0]    reg_weight_3_39;
wire signed[31:0]    reg_psum_3_39;
wire signed[31:0]    reg_weight_3_40;
wire signed[31:0]    reg_psum_3_40;
wire signed[31:0]    reg_weight_3_41;
wire signed[31:0]    reg_psum_3_41;
wire signed[31:0]    reg_weight_3_42;
wire signed[31:0]    reg_psum_3_42;
wire signed[31:0]    reg_weight_3_43;
wire signed[31:0]    reg_psum_3_43;
wire signed[31:0]    reg_weight_3_44;
wire signed[31:0]    reg_psum_3_44;
wire signed[31:0]    reg_weight_3_45;
wire signed[31:0]    reg_psum_3_45;
wire signed[31:0]    reg_weight_3_46;
wire signed[31:0]    reg_psum_3_46;
wire signed[31:0]    reg_weight_3_47;
wire signed[31:0]    reg_psum_3_47;
wire signed[31:0]    reg_weight_3_48;
wire signed[31:0]    reg_psum_3_48;
wire signed[31:0]    reg_weight_3_49;
wire signed[31:0]    reg_psum_3_49;
wire signed[31:0]    reg_weight_3_50;
wire signed[31:0]    reg_psum_3_50;
wire signed[31:0]    reg_weight_3_51;
wire signed[31:0]    reg_psum_3_51;
wire signed[31:0]    reg_weight_3_52;
wire signed[31:0]    reg_psum_3_52;
wire signed[31:0]    reg_weight_3_53;
wire signed[31:0]    reg_psum_3_53;
wire signed[31:0]    reg_weight_3_54;
wire signed[31:0]    reg_psum_3_54;
wire signed[31:0]    reg_weight_3_55;
wire signed[31:0]    reg_psum_3_55;
wire signed[31:0]    reg_weight_3_56;
wire signed[31:0]    reg_psum_3_56;
wire signed[31:0]    reg_weight_3_57;
wire signed[31:0]    reg_psum_3_57;
wire signed[31:0]    reg_weight_3_58;
wire signed[31:0]    reg_psum_3_58;
wire signed[31:0]    reg_weight_3_59;
wire signed[31:0]    reg_psum_3_59;
wire signed[31:0]    reg_weight_3_60;
wire signed[31:0]    reg_psum_3_60;
wire signed[31:0]    reg_weight_3_61;
wire signed[31:0]    reg_psum_3_61;
wire signed[31:0]    reg_weight_3_62;
wire signed[31:0]    reg_psum_3_62;
wire signed[31:0]    reg_weight_3_63;
wire signed[31:0]    reg_psum_3_63;
wire signed[31:0]    reg_weight_4_0;
wire signed[31:0]    reg_psum_4_0;
wire signed[31:0]    reg_weight_4_1;
wire signed[31:0]    reg_psum_4_1;
wire signed[31:0]    reg_weight_4_2;
wire signed[31:0]    reg_psum_4_2;
wire signed[31:0]    reg_weight_4_3;
wire signed[31:0]    reg_psum_4_3;
wire signed[31:0]    reg_weight_4_4;
wire signed[31:0]    reg_psum_4_4;
wire signed[31:0]    reg_weight_4_5;
wire signed[31:0]    reg_psum_4_5;
wire signed[31:0]    reg_weight_4_6;
wire signed[31:0]    reg_psum_4_6;
wire signed[31:0]    reg_weight_4_7;
wire signed[31:0]    reg_psum_4_7;
wire signed[31:0]    reg_weight_4_8;
wire signed[31:0]    reg_psum_4_8;
wire signed[31:0]    reg_weight_4_9;
wire signed[31:0]    reg_psum_4_9;
wire signed[31:0]    reg_weight_4_10;
wire signed[31:0]    reg_psum_4_10;
wire signed[31:0]    reg_weight_4_11;
wire signed[31:0]    reg_psum_4_11;
wire signed[31:0]    reg_weight_4_12;
wire signed[31:0]    reg_psum_4_12;
wire signed[31:0]    reg_weight_4_13;
wire signed[31:0]    reg_psum_4_13;
wire signed[31:0]    reg_weight_4_14;
wire signed[31:0]    reg_psum_4_14;
wire signed[31:0]    reg_weight_4_15;
wire signed[31:0]    reg_psum_4_15;
wire signed[31:0]    reg_weight_4_16;
wire signed[31:0]    reg_psum_4_16;
wire signed[31:0]    reg_weight_4_17;
wire signed[31:0]    reg_psum_4_17;
wire signed[31:0]    reg_weight_4_18;
wire signed[31:0]    reg_psum_4_18;
wire signed[31:0]    reg_weight_4_19;
wire signed[31:0]    reg_psum_4_19;
wire signed[31:0]    reg_weight_4_20;
wire signed[31:0]    reg_psum_4_20;
wire signed[31:0]    reg_weight_4_21;
wire signed[31:0]    reg_psum_4_21;
wire signed[31:0]    reg_weight_4_22;
wire signed[31:0]    reg_psum_4_22;
wire signed[31:0]    reg_weight_4_23;
wire signed[31:0]    reg_psum_4_23;
wire signed[31:0]    reg_weight_4_24;
wire signed[31:0]    reg_psum_4_24;
wire signed[31:0]    reg_weight_4_25;
wire signed[31:0]    reg_psum_4_25;
wire signed[31:0]    reg_weight_4_26;
wire signed[31:0]    reg_psum_4_26;
wire signed[31:0]    reg_weight_4_27;
wire signed[31:0]    reg_psum_4_27;
wire signed[31:0]    reg_weight_4_28;
wire signed[31:0]    reg_psum_4_28;
wire signed[31:0]    reg_weight_4_29;
wire signed[31:0]    reg_psum_4_29;
wire signed[31:0]    reg_weight_4_30;
wire signed[31:0]    reg_psum_4_30;
wire signed[31:0]    reg_weight_4_31;
wire signed[31:0]    reg_psum_4_31;
wire signed[31:0]    reg_weight_4_32;
wire signed[31:0]    reg_psum_4_32;
wire signed[31:0]    reg_weight_4_33;
wire signed[31:0]    reg_psum_4_33;
wire signed[31:0]    reg_weight_4_34;
wire signed[31:0]    reg_psum_4_34;
wire signed[31:0]    reg_weight_4_35;
wire signed[31:0]    reg_psum_4_35;
wire signed[31:0]    reg_weight_4_36;
wire signed[31:0]    reg_psum_4_36;
wire signed[31:0]    reg_weight_4_37;
wire signed[31:0]    reg_psum_4_37;
wire signed[31:0]    reg_weight_4_38;
wire signed[31:0]    reg_psum_4_38;
wire signed[31:0]    reg_weight_4_39;
wire signed[31:0]    reg_psum_4_39;
wire signed[31:0]    reg_weight_4_40;
wire signed[31:0]    reg_psum_4_40;
wire signed[31:0]    reg_weight_4_41;
wire signed[31:0]    reg_psum_4_41;
wire signed[31:0]    reg_weight_4_42;
wire signed[31:0]    reg_psum_4_42;
wire signed[31:0]    reg_weight_4_43;
wire signed[31:0]    reg_psum_4_43;
wire signed[31:0]    reg_weight_4_44;
wire signed[31:0]    reg_psum_4_44;
wire signed[31:0]    reg_weight_4_45;
wire signed[31:0]    reg_psum_4_45;
wire signed[31:0]    reg_weight_4_46;
wire signed[31:0]    reg_psum_4_46;
wire signed[31:0]    reg_weight_4_47;
wire signed[31:0]    reg_psum_4_47;
wire signed[31:0]    reg_weight_4_48;
wire signed[31:0]    reg_psum_4_48;
wire signed[31:0]    reg_weight_4_49;
wire signed[31:0]    reg_psum_4_49;
wire signed[31:0]    reg_weight_4_50;
wire signed[31:0]    reg_psum_4_50;
wire signed[31:0]    reg_weight_4_51;
wire signed[31:0]    reg_psum_4_51;
wire signed[31:0]    reg_weight_4_52;
wire signed[31:0]    reg_psum_4_52;
wire signed[31:0]    reg_weight_4_53;
wire signed[31:0]    reg_psum_4_53;
wire signed[31:0]    reg_weight_4_54;
wire signed[31:0]    reg_psum_4_54;
wire signed[31:0]    reg_weight_4_55;
wire signed[31:0]    reg_psum_4_55;
wire signed[31:0]    reg_weight_4_56;
wire signed[31:0]    reg_psum_4_56;
wire signed[31:0]    reg_weight_4_57;
wire signed[31:0]    reg_psum_4_57;
wire signed[31:0]    reg_weight_4_58;
wire signed[31:0]    reg_psum_4_58;
wire signed[31:0]    reg_weight_4_59;
wire signed[31:0]    reg_psum_4_59;
wire signed[31:0]    reg_weight_4_60;
wire signed[31:0]    reg_psum_4_60;
wire signed[31:0]    reg_weight_4_61;
wire signed[31:0]    reg_psum_4_61;
wire signed[31:0]    reg_weight_4_62;
wire signed[31:0]    reg_psum_4_62;
wire signed[31:0]    reg_weight_4_63;
wire signed[31:0]    reg_psum_4_63;
wire signed[31:0]    reg_weight_5_0;
wire signed[31:0]    reg_psum_5_0;
wire signed[31:0]    reg_weight_5_1;
wire signed[31:0]    reg_psum_5_1;
wire signed[31:0]    reg_weight_5_2;
wire signed[31:0]    reg_psum_5_2;
wire signed[31:0]    reg_weight_5_3;
wire signed[31:0]    reg_psum_5_3;
wire signed[31:0]    reg_weight_5_4;
wire signed[31:0]    reg_psum_5_4;
wire signed[31:0]    reg_weight_5_5;
wire signed[31:0]    reg_psum_5_5;
wire signed[31:0]    reg_weight_5_6;
wire signed[31:0]    reg_psum_5_6;
wire signed[31:0]    reg_weight_5_7;
wire signed[31:0]    reg_psum_5_7;
wire signed[31:0]    reg_weight_5_8;
wire signed[31:0]    reg_psum_5_8;
wire signed[31:0]    reg_weight_5_9;
wire signed[31:0]    reg_psum_5_9;
wire signed[31:0]    reg_weight_5_10;
wire signed[31:0]    reg_psum_5_10;
wire signed[31:0]    reg_weight_5_11;
wire signed[31:0]    reg_psum_5_11;
wire signed[31:0]    reg_weight_5_12;
wire signed[31:0]    reg_psum_5_12;
wire signed[31:0]    reg_weight_5_13;
wire signed[31:0]    reg_psum_5_13;
wire signed[31:0]    reg_weight_5_14;
wire signed[31:0]    reg_psum_5_14;
wire signed[31:0]    reg_weight_5_15;
wire signed[31:0]    reg_psum_5_15;
wire signed[31:0]    reg_weight_5_16;
wire signed[31:0]    reg_psum_5_16;
wire signed[31:0]    reg_weight_5_17;
wire signed[31:0]    reg_psum_5_17;
wire signed[31:0]    reg_weight_5_18;
wire signed[31:0]    reg_psum_5_18;
wire signed[31:0]    reg_weight_5_19;
wire signed[31:0]    reg_psum_5_19;
wire signed[31:0]    reg_weight_5_20;
wire signed[31:0]    reg_psum_5_20;
wire signed[31:0]    reg_weight_5_21;
wire signed[31:0]    reg_psum_5_21;
wire signed[31:0]    reg_weight_5_22;
wire signed[31:0]    reg_psum_5_22;
wire signed[31:0]    reg_weight_5_23;
wire signed[31:0]    reg_psum_5_23;
wire signed[31:0]    reg_weight_5_24;
wire signed[31:0]    reg_psum_5_24;
wire signed[31:0]    reg_weight_5_25;
wire signed[31:0]    reg_psum_5_25;
wire signed[31:0]    reg_weight_5_26;
wire signed[31:0]    reg_psum_5_26;
wire signed[31:0]    reg_weight_5_27;
wire signed[31:0]    reg_psum_5_27;
wire signed[31:0]    reg_weight_5_28;
wire signed[31:0]    reg_psum_5_28;
wire signed[31:0]    reg_weight_5_29;
wire signed[31:0]    reg_psum_5_29;
wire signed[31:0]    reg_weight_5_30;
wire signed[31:0]    reg_psum_5_30;
wire signed[31:0]    reg_weight_5_31;
wire signed[31:0]    reg_psum_5_31;
wire signed[31:0]    reg_weight_5_32;
wire signed[31:0]    reg_psum_5_32;
wire signed[31:0]    reg_weight_5_33;
wire signed[31:0]    reg_psum_5_33;
wire signed[31:0]    reg_weight_5_34;
wire signed[31:0]    reg_psum_5_34;
wire signed[31:0]    reg_weight_5_35;
wire signed[31:0]    reg_psum_5_35;
wire signed[31:0]    reg_weight_5_36;
wire signed[31:0]    reg_psum_5_36;
wire signed[31:0]    reg_weight_5_37;
wire signed[31:0]    reg_psum_5_37;
wire signed[31:0]    reg_weight_5_38;
wire signed[31:0]    reg_psum_5_38;
wire signed[31:0]    reg_weight_5_39;
wire signed[31:0]    reg_psum_5_39;
wire signed[31:0]    reg_weight_5_40;
wire signed[31:0]    reg_psum_5_40;
wire signed[31:0]    reg_weight_5_41;
wire signed[31:0]    reg_psum_5_41;
wire signed[31:0]    reg_weight_5_42;
wire signed[31:0]    reg_psum_5_42;
wire signed[31:0]    reg_weight_5_43;
wire signed[31:0]    reg_psum_5_43;
wire signed[31:0]    reg_weight_5_44;
wire signed[31:0]    reg_psum_5_44;
wire signed[31:0]    reg_weight_5_45;
wire signed[31:0]    reg_psum_5_45;
wire signed[31:0]    reg_weight_5_46;
wire signed[31:0]    reg_psum_5_46;
wire signed[31:0]    reg_weight_5_47;
wire signed[31:0]    reg_psum_5_47;
wire signed[31:0]    reg_weight_5_48;
wire signed[31:0]    reg_psum_5_48;
wire signed[31:0]    reg_weight_5_49;
wire signed[31:0]    reg_psum_5_49;
wire signed[31:0]    reg_weight_5_50;
wire signed[31:0]    reg_psum_5_50;
wire signed[31:0]    reg_weight_5_51;
wire signed[31:0]    reg_psum_5_51;
wire signed[31:0]    reg_weight_5_52;
wire signed[31:0]    reg_psum_5_52;
wire signed[31:0]    reg_weight_5_53;
wire signed[31:0]    reg_psum_5_53;
wire signed[31:0]    reg_weight_5_54;
wire signed[31:0]    reg_psum_5_54;
wire signed[31:0]    reg_weight_5_55;
wire signed[31:0]    reg_psum_5_55;
wire signed[31:0]    reg_weight_5_56;
wire signed[31:0]    reg_psum_5_56;
wire signed[31:0]    reg_weight_5_57;
wire signed[31:0]    reg_psum_5_57;
wire signed[31:0]    reg_weight_5_58;
wire signed[31:0]    reg_psum_5_58;
wire signed[31:0]    reg_weight_5_59;
wire signed[31:0]    reg_psum_5_59;
wire signed[31:0]    reg_weight_5_60;
wire signed[31:0]    reg_psum_5_60;
wire signed[31:0]    reg_weight_5_61;
wire signed[31:0]    reg_psum_5_61;
wire signed[31:0]    reg_weight_5_62;
wire signed[31:0]    reg_psum_5_62;
wire signed[31:0]    reg_weight_5_63;
wire signed[31:0]    reg_psum_5_63;
wire signed[31:0]    reg_weight_6_0;
wire signed[31:0]    reg_psum_6_0;
wire signed[31:0]    reg_weight_6_1;
wire signed[31:0]    reg_psum_6_1;
wire signed[31:0]    reg_weight_6_2;
wire signed[31:0]    reg_psum_6_2;
wire signed[31:0]    reg_weight_6_3;
wire signed[31:0]    reg_psum_6_3;
wire signed[31:0]    reg_weight_6_4;
wire signed[31:0]    reg_psum_6_4;
wire signed[31:0]    reg_weight_6_5;
wire signed[31:0]    reg_psum_6_5;
wire signed[31:0]    reg_weight_6_6;
wire signed[31:0]    reg_psum_6_6;
wire signed[31:0]    reg_weight_6_7;
wire signed[31:0]    reg_psum_6_7;
wire signed[31:0]    reg_weight_6_8;
wire signed[31:0]    reg_psum_6_8;
wire signed[31:0]    reg_weight_6_9;
wire signed[31:0]    reg_psum_6_9;
wire signed[31:0]    reg_weight_6_10;
wire signed[31:0]    reg_psum_6_10;
wire signed[31:0]    reg_weight_6_11;
wire signed[31:0]    reg_psum_6_11;
wire signed[31:0]    reg_weight_6_12;
wire signed[31:0]    reg_psum_6_12;
wire signed[31:0]    reg_weight_6_13;
wire signed[31:0]    reg_psum_6_13;
wire signed[31:0]    reg_weight_6_14;
wire signed[31:0]    reg_psum_6_14;
wire signed[31:0]    reg_weight_6_15;
wire signed[31:0]    reg_psum_6_15;
wire signed[31:0]    reg_weight_6_16;
wire signed[31:0]    reg_psum_6_16;
wire signed[31:0]    reg_weight_6_17;
wire signed[31:0]    reg_psum_6_17;
wire signed[31:0]    reg_weight_6_18;
wire signed[31:0]    reg_psum_6_18;
wire signed[31:0]    reg_weight_6_19;
wire signed[31:0]    reg_psum_6_19;
wire signed[31:0]    reg_weight_6_20;
wire signed[31:0]    reg_psum_6_20;
wire signed[31:0]    reg_weight_6_21;
wire signed[31:0]    reg_psum_6_21;
wire signed[31:0]    reg_weight_6_22;
wire signed[31:0]    reg_psum_6_22;
wire signed[31:0]    reg_weight_6_23;
wire signed[31:0]    reg_psum_6_23;
wire signed[31:0]    reg_weight_6_24;
wire signed[31:0]    reg_psum_6_24;
wire signed[31:0]    reg_weight_6_25;
wire signed[31:0]    reg_psum_6_25;
wire signed[31:0]    reg_weight_6_26;
wire signed[31:0]    reg_psum_6_26;
wire signed[31:0]    reg_weight_6_27;
wire signed[31:0]    reg_psum_6_27;
wire signed[31:0]    reg_weight_6_28;
wire signed[31:0]    reg_psum_6_28;
wire signed[31:0]    reg_weight_6_29;
wire signed[31:0]    reg_psum_6_29;
wire signed[31:0]    reg_weight_6_30;
wire signed[31:0]    reg_psum_6_30;
wire signed[31:0]    reg_weight_6_31;
wire signed[31:0]    reg_psum_6_31;
wire signed[31:0]    reg_weight_6_32;
wire signed[31:0]    reg_psum_6_32;
wire signed[31:0]    reg_weight_6_33;
wire signed[31:0]    reg_psum_6_33;
wire signed[31:0]    reg_weight_6_34;
wire signed[31:0]    reg_psum_6_34;
wire signed[31:0]    reg_weight_6_35;
wire signed[31:0]    reg_psum_6_35;
wire signed[31:0]    reg_weight_6_36;
wire signed[31:0]    reg_psum_6_36;
wire signed[31:0]    reg_weight_6_37;
wire signed[31:0]    reg_psum_6_37;
wire signed[31:0]    reg_weight_6_38;
wire signed[31:0]    reg_psum_6_38;
wire signed[31:0]    reg_weight_6_39;
wire signed[31:0]    reg_psum_6_39;
wire signed[31:0]    reg_weight_6_40;
wire signed[31:0]    reg_psum_6_40;
wire signed[31:0]    reg_weight_6_41;
wire signed[31:0]    reg_psum_6_41;
wire signed[31:0]    reg_weight_6_42;
wire signed[31:0]    reg_psum_6_42;
wire signed[31:0]    reg_weight_6_43;
wire signed[31:0]    reg_psum_6_43;
wire signed[31:0]    reg_weight_6_44;
wire signed[31:0]    reg_psum_6_44;
wire signed[31:0]    reg_weight_6_45;
wire signed[31:0]    reg_psum_6_45;
wire signed[31:0]    reg_weight_6_46;
wire signed[31:0]    reg_psum_6_46;
wire signed[31:0]    reg_weight_6_47;
wire signed[31:0]    reg_psum_6_47;
wire signed[31:0]    reg_weight_6_48;
wire signed[31:0]    reg_psum_6_48;
wire signed[31:0]    reg_weight_6_49;
wire signed[31:0]    reg_psum_6_49;
wire signed[31:0]    reg_weight_6_50;
wire signed[31:0]    reg_psum_6_50;
wire signed[31:0]    reg_weight_6_51;
wire signed[31:0]    reg_psum_6_51;
wire signed[31:0]    reg_weight_6_52;
wire signed[31:0]    reg_psum_6_52;
wire signed[31:0]    reg_weight_6_53;
wire signed[31:0]    reg_psum_6_53;
wire signed[31:0]    reg_weight_6_54;
wire signed[31:0]    reg_psum_6_54;
wire signed[31:0]    reg_weight_6_55;
wire signed[31:0]    reg_psum_6_55;
wire signed[31:0]    reg_weight_6_56;
wire signed[31:0]    reg_psum_6_56;
wire signed[31:0]    reg_weight_6_57;
wire signed[31:0]    reg_psum_6_57;
wire signed[31:0]    reg_weight_6_58;
wire signed[31:0]    reg_psum_6_58;
wire signed[31:0]    reg_weight_6_59;
wire signed[31:0]    reg_psum_6_59;
wire signed[31:0]    reg_weight_6_60;
wire signed[31:0]    reg_psum_6_60;
wire signed[31:0]    reg_weight_6_61;
wire signed[31:0]    reg_psum_6_61;
wire signed[31:0]    reg_weight_6_62;
wire signed[31:0]    reg_psum_6_62;
wire signed[31:0]    reg_weight_6_63;
wire signed[31:0]    reg_psum_6_63;
wire signed[31:0]    reg_weight_7_0;
wire signed[31:0]    reg_psum_7_0;
wire signed[31:0]    reg_weight_7_1;
wire signed[31:0]    reg_psum_7_1;
wire signed[31:0]    reg_weight_7_2;
wire signed[31:0]    reg_psum_7_2;
wire signed[31:0]    reg_weight_7_3;
wire signed[31:0]    reg_psum_7_3;
wire signed[31:0]    reg_weight_7_4;
wire signed[31:0]    reg_psum_7_4;
wire signed[31:0]    reg_weight_7_5;
wire signed[31:0]    reg_psum_7_5;
wire signed[31:0]    reg_weight_7_6;
wire signed[31:0]    reg_psum_7_6;
wire signed[31:0]    reg_weight_7_7;
wire signed[31:0]    reg_psum_7_7;
wire signed[31:0]    reg_weight_7_8;
wire signed[31:0]    reg_psum_7_8;
wire signed[31:0]    reg_weight_7_9;
wire signed[31:0]    reg_psum_7_9;
wire signed[31:0]    reg_weight_7_10;
wire signed[31:0]    reg_psum_7_10;
wire signed[31:0]    reg_weight_7_11;
wire signed[31:0]    reg_psum_7_11;
wire signed[31:0]    reg_weight_7_12;
wire signed[31:0]    reg_psum_7_12;
wire signed[31:0]    reg_weight_7_13;
wire signed[31:0]    reg_psum_7_13;
wire signed[31:0]    reg_weight_7_14;
wire signed[31:0]    reg_psum_7_14;
wire signed[31:0]    reg_weight_7_15;
wire signed[31:0]    reg_psum_7_15;
wire signed[31:0]    reg_weight_7_16;
wire signed[31:0]    reg_psum_7_16;
wire signed[31:0]    reg_weight_7_17;
wire signed[31:0]    reg_psum_7_17;
wire signed[31:0]    reg_weight_7_18;
wire signed[31:0]    reg_psum_7_18;
wire signed[31:0]    reg_weight_7_19;
wire signed[31:0]    reg_psum_7_19;
wire signed[31:0]    reg_weight_7_20;
wire signed[31:0]    reg_psum_7_20;
wire signed[31:0]    reg_weight_7_21;
wire signed[31:0]    reg_psum_7_21;
wire signed[31:0]    reg_weight_7_22;
wire signed[31:0]    reg_psum_7_22;
wire signed[31:0]    reg_weight_7_23;
wire signed[31:0]    reg_psum_7_23;
wire signed[31:0]    reg_weight_7_24;
wire signed[31:0]    reg_psum_7_24;
wire signed[31:0]    reg_weight_7_25;
wire signed[31:0]    reg_psum_7_25;
wire signed[31:0]    reg_weight_7_26;
wire signed[31:0]    reg_psum_7_26;
wire signed[31:0]    reg_weight_7_27;
wire signed[31:0]    reg_psum_7_27;
wire signed[31:0]    reg_weight_7_28;
wire signed[31:0]    reg_psum_7_28;
wire signed[31:0]    reg_weight_7_29;
wire signed[31:0]    reg_psum_7_29;
wire signed[31:0]    reg_weight_7_30;
wire signed[31:0]    reg_psum_7_30;
wire signed[31:0]    reg_weight_7_31;
wire signed[31:0]    reg_psum_7_31;
wire signed[31:0]    reg_weight_7_32;
wire signed[31:0]    reg_psum_7_32;
wire signed[31:0]    reg_weight_7_33;
wire signed[31:0]    reg_psum_7_33;
wire signed[31:0]    reg_weight_7_34;
wire signed[31:0]    reg_psum_7_34;
wire signed[31:0]    reg_weight_7_35;
wire signed[31:0]    reg_psum_7_35;
wire signed[31:0]    reg_weight_7_36;
wire signed[31:0]    reg_psum_7_36;
wire signed[31:0]    reg_weight_7_37;
wire signed[31:0]    reg_psum_7_37;
wire signed[31:0]    reg_weight_7_38;
wire signed[31:0]    reg_psum_7_38;
wire signed[31:0]    reg_weight_7_39;
wire signed[31:0]    reg_psum_7_39;
wire signed[31:0]    reg_weight_7_40;
wire signed[31:0]    reg_psum_7_40;
wire signed[31:0]    reg_weight_7_41;
wire signed[31:0]    reg_psum_7_41;
wire signed[31:0]    reg_weight_7_42;
wire signed[31:0]    reg_psum_7_42;
wire signed[31:0]    reg_weight_7_43;
wire signed[31:0]    reg_psum_7_43;
wire signed[31:0]    reg_weight_7_44;
wire signed[31:0]    reg_psum_7_44;
wire signed[31:0]    reg_weight_7_45;
wire signed[31:0]    reg_psum_7_45;
wire signed[31:0]    reg_weight_7_46;
wire signed[31:0]    reg_psum_7_46;
wire signed[31:0]    reg_weight_7_47;
wire signed[31:0]    reg_psum_7_47;
wire signed[31:0]    reg_weight_7_48;
wire signed[31:0]    reg_psum_7_48;
wire signed[31:0]    reg_weight_7_49;
wire signed[31:0]    reg_psum_7_49;
wire signed[31:0]    reg_weight_7_50;
wire signed[31:0]    reg_psum_7_50;
wire signed[31:0]    reg_weight_7_51;
wire signed[31:0]    reg_psum_7_51;
wire signed[31:0]    reg_weight_7_52;
wire signed[31:0]    reg_psum_7_52;
wire signed[31:0]    reg_weight_7_53;
wire signed[31:0]    reg_psum_7_53;
wire signed[31:0]    reg_weight_7_54;
wire signed[31:0]    reg_psum_7_54;
wire signed[31:0]    reg_weight_7_55;
wire signed[31:0]    reg_psum_7_55;
wire signed[31:0]    reg_weight_7_56;
wire signed[31:0]    reg_psum_7_56;
wire signed[31:0]    reg_weight_7_57;
wire signed[31:0]    reg_psum_7_57;
wire signed[31:0]    reg_weight_7_58;
wire signed[31:0]    reg_psum_7_58;
wire signed[31:0]    reg_weight_7_59;
wire signed[31:0]    reg_psum_7_59;
wire signed[31:0]    reg_weight_7_60;
wire signed[31:0]    reg_psum_7_60;
wire signed[31:0]    reg_weight_7_61;
wire signed[31:0]    reg_psum_7_61;
wire signed[31:0]    reg_weight_7_62;
wire signed[31:0]    reg_psum_7_62;
wire signed[31:0]    reg_weight_7_63;
wire signed[31:0]    reg_psum_7_63;
wire signed[31:0]    reg_weight_8_0;
wire signed[31:0]    reg_psum_8_0;
wire signed[31:0]    reg_weight_8_1;
wire signed[31:0]    reg_psum_8_1;
wire signed[31:0]    reg_weight_8_2;
wire signed[31:0]    reg_psum_8_2;
wire signed[31:0]    reg_weight_8_3;
wire signed[31:0]    reg_psum_8_3;
wire signed[31:0]    reg_weight_8_4;
wire signed[31:0]    reg_psum_8_4;
wire signed[31:0]    reg_weight_8_5;
wire signed[31:0]    reg_psum_8_5;
wire signed[31:0]    reg_weight_8_6;
wire signed[31:0]    reg_psum_8_6;
wire signed[31:0]    reg_weight_8_7;
wire signed[31:0]    reg_psum_8_7;
wire signed[31:0]    reg_weight_8_8;
wire signed[31:0]    reg_psum_8_8;
wire signed[31:0]    reg_weight_8_9;
wire signed[31:0]    reg_psum_8_9;
wire signed[31:0]    reg_weight_8_10;
wire signed[31:0]    reg_psum_8_10;
wire signed[31:0]    reg_weight_8_11;
wire signed[31:0]    reg_psum_8_11;
wire signed[31:0]    reg_weight_8_12;
wire signed[31:0]    reg_psum_8_12;
wire signed[31:0]    reg_weight_8_13;
wire signed[31:0]    reg_psum_8_13;
wire signed[31:0]    reg_weight_8_14;
wire signed[31:0]    reg_psum_8_14;
wire signed[31:0]    reg_weight_8_15;
wire signed[31:0]    reg_psum_8_15;
wire signed[31:0]    reg_weight_8_16;
wire signed[31:0]    reg_psum_8_16;
wire signed[31:0]    reg_weight_8_17;
wire signed[31:0]    reg_psum_8_17;
wire signed[31:0]    reg_weight_8_18;
wire signed[31:0]    reg_psum_8_18;
wire signed[31:0]    reg_weight_8_19;
wire signed[31:0]    reg_psum_8_19;
wire signed[31:0]    reg_weight_8_20;
wire signed[31:0]    reg_psum_8_20;
wire signed[31:0]    reg_weight_8_21;
wire signed[31:0]    reg_psum_8_21;
wire signed[31:0]    reg_weight_8_22;
wire signed[31:0]    reg_psum_8_22;
wire signed[31:0]    reg_weight_8_23;
wire signed[31:0]    reg_psum_8_23;
wire signed[31:0]    reg_weight_8_24;
wire signed[31:0]    reg_psum_8_24;
wire signed[31:0]    reg_weight_8_25;
wire signed[31:0]    reg_psum_8_25;
wire signed[31:0]    reg_weight_8_26;
wire signed[31:0]    reg_psum_8_26;
wire signed[31:0]    reg_weight_8_27;
wire signed[31:0]    reg_psum_8_27;
wire signed[31:0]    reg_weight_8_28;
wire signed[31:0]    reg_psum_8_28;
wire signed[31:0]    reg_weight_8_29;
wire signed[31:0]    reg_psum_8_29;
wire signed[31:0]    reg_weight_8_30;
wire signed[31:0]    reg_psum_8_30;
wire signed[31:0]    reg_weight_8_31;
wire signed[31:0]    reg_psum_8_31;
wire signed[31:0]    reg_weight_8_32;
wire signed[31:0]    reg_psum_8_32;
wire signed[31:0]    reg_weight_8_33;
wire signed[31:0]    reg_psum_8_33;
wire signed[31:0]    reg_weight_8_34;
wire signed[31:0]    reg_psum_8_34;
wire signed[31:0]    reg_weight_8_35;
wire signed[31:0]    reg_psum_8_35;
wire signed[31:0]    reg_weight_8_36;
wire signed[31:0]    reg_psum_8_36;
wire signed[31:0]    reg_weight_8_37;
wire signed[31:0]    reg_psum_8_37;
wire signed[31:0]    reg_weight_8_38;
wire signed[31:0]    reg_psum_8_38;
wire signed[31:0]    reg_weight_8_39;
wire signed[31:0]    reg_psum_8_39;
wire signed[31:0]    reg_weight_8_40;
wire signed[31:0]    reg_psum_8_40;
wire signed[31:0]    reg_weight_8_41;
wire signed[31:0]    reg_psum_8_41;
wire signed[31:0]    reg_weight_8_42;
wire signed[31:0]    reg_psum_8_42;
wire signed[31:0]    reg_weight_8_43;
wire signed[31:0]    reg_psum_8_43;
wire signed[31:0]    reg_weight_8_44;
wire signed[31:0]    reg_psum_8_44;
wire signed[31:0]    reg_weight_8_45;
wire signed[31:0]    reg_psum_8_45;
wire signed[31:0]    reg_weight_8_46;
wire signed[31:0]    reg_psum_8_46;
wire signed[31:0]    reg_weight_8_47;
wire signed[31:0]    reg_psum_8_47;
wire signed[31:0]    reg_weight_8_48;
wire signed[31:0]    reg_psum_8_48;
wire signed[31:0]    reg_weight_8_49;
wire signed[31:0]    reg_psum_8_49;
wire signed[31:0]    reg_weight_8_50;
wire signed[31:0]    reg_psum_8_50;
wire signed[31:0]    reg_weight_8_51;
wire signed[31:0]    reg_psum_8_51;
wire signed[31:0]    reg_weight_8_52;
wire signed[31:0]    reg_psum_8_52;
wire signed[31:0]    reg_weight_8_53;
wire signed[31:0]    reg_psum_8_53;
wire signed[31:0]    reg_weight_8_54;
wire signed[31:0]    reg_psum_8_54;
wire signed[31:0]    reg_weight_8_55;
wire signed[31:0]    reg_psum_8_55;
wire signed[31:0]    reg_weight_8_56;
wire signed[31:0]    reg_psum_8_56;
wire signed[31:0]    reg_weight_8_57;
wire signed[31:0]    reg_psum_8_57;
wire signed[31:0]    reg_weight_8_58;
wire signed[31:0]    reg_psum_8_58;
wire signed[31:0]    reg_weight_8_59;
wire signed[31:0]    reg_psum_8_59;
wire signed[31:0]    reg_weight_8_60;
wire signed[31:0]    reg_psum_8_60;
wire signed[31:0]    reg_weight_8_61;
wire signed[31:0]    reg_psum_8_61;
wire signed[31:0]    reg_weight_8_62;
wire signed[31:0]    reg_psum_8_62;
wire signed[31:0]    reg_weight_8_63;
wire signed[31:0]    reg_psum_8_63;
wire signed[31:0]    reg_weight_9_0;
wire signed[31:0]    reg_psum_9_0;
wire signed[31:0]    reg_weight_9_1;
wire signed[31:0]    reg_psum_9_1;
wire signed[31:0]    reg_weight_9_2;
wire signed[31:0]    reg_psum_9_2;
wire signed[31:0]    reg_weight_9_3;
wire signed[31:0]    reg_psum_9_3;
wire signed[31:0]    reg_weight_9_4;
wire signed[31:0]    reg_psum_9_4;
wire signed[31:0]    reg_weight_9_5;
wire signed[31:0]    reg_psum_9_5;
wire signed[31:0]    reg_weight_9_6;
wire signed[31:0]    reg_psum_9_6;
wire signed[31:0]    reg_weight_9_7;
wire signed[31:0]    reg_psum_9_7;
wire signed[31:0]    reg_weight_9_8;
wire signed[31:0]    reg_psum_9_8;
wire signed[31:0]    reg_weight_9_9;
wire signed[31:0]    reg_psum_9_9;
wire signed[31:0]    reg_weight_9_10;
wire signed[31:0]    reg_psum_9_10;
wire signed[31:0]    reg_weight_9_11;
wire signed[31:0]    reg_psum_9_11;
wire signed[31:0]    reg_weight_9_12;
wire signed[31:0]    reg_psum_9_12;
wire signed[31:0]    reg_weight_9_13;
wire signed[31:0]    reg_psum_9_13;
wire signed[31:0]    reg_weight_9_14;
wire signed[31:0]    reg_psum_9_14;
wire signed[31:0]    reg_weight_9_15;
wire signed[31:0]    reg_psum_9_15;
wire signed[31:0]    reg_weight_9_16;
wire signed[31:0]    reg_psum_9_16;
wire signed[31:0]    reg_weight_9_17;
wire signed[31:0]    reg_psum_9_17;
wire signed[31:0]    reg_weight_9_18;
wire signed[31:0]    reg_psum_9_18;
wire signed[31:0]    reg_weight_9_19;
wire signed[31:0]    reg_psum_9_19;
wire signed[31:0]    reg_weight_9_20;
wire signed[31:0]    reg_psum_9_20;
wire signed[31:0]    reg_weight_9_21;
wire signed[31:0]    reg_psum_9_21;
wire signed[31:0]    reg_weight_9_22;
wire signed[31:0]    reg_psum_9_22;
wire signed[31:0]    reg_weight_9_23;
wire signed[31:0]    reg_psum_9_23;
wire signed[31:0]    reg_weight_9_24;
wire signed[31:0]    reg_psum_9_24;
wire signed[31:0]    reg_weight_9_25;
wire signed[31:0]    reg_psum_9_25;
wire signed[31:0]    reg_weight_9_26;
wire signed[31:0]    reg_psum_9_26;
wire signed[31:0]    reg_weight_9_27;
wire signed[31:0]    reg_psum_9_27;
wire signed[31:0]    reg_weight_9_28;
wire signed[31:0]    reg_psum_9_28;
wire signed[31:0]    reg_weight_9_29;
wire signed[31:0]    reg_psum_9_29;
wire signed[31:0]    reg_weight_9_30;
wire signed[31:0]    reg_psum_9_30;
wire signed[31:0]    reg_weight_9_31;
wire signed[31:0]    reg_psum_9_31;
wire signed[31:0]    reg_weight_9_32;
wire signed[31:0]    reg_psum_9_32;
wire signed[31:0]    reg_weight_9_33;
wire signed[31:0]    reg_psum_9_33;
wire signed[31:0]    reg_weight_9_34;
wire signed[31:0]    reg_psum_9_34;
wire signed[31:0]    reg_weight_9_35;
wire signed[31:0]    reg_psum_9_35;
wire signed[31:0]    reg_weight_9_36;
wire signed[31:0]    reg_psum_9_36;
wire signed[31:0]    reg_weight_9_37;
wire signed[31:0]    reg_psum_9_37;
wire signed[31:0]    reg_weight_9_38;
wire signed[31:0]    reg_psum_9_38;
wire signed[31:0]    reg_weight_9_39;
wire signed[31:0]    reg_psum_9_39;
wire signed[31:0]    reg_weight_9_40;
wire signed[31:0]    reg_psum_9_40;
wire signed[31:0]    reg_weight_9_41;
wire signed[31:0]    reg_psum_9_41;
wire signed[31:0]    reg_weight_9_42;
wire signed[31:0]    reg_psum_9_42;
wire signed[31:0]    reg_weight_9_43;
wire signed[31:0]    reg_psum_9_43;
wire signed[31:0]    reg_weight_9_44;
wire signed[31:0]    reg_psum_9_44;
wire signed[31:0]    reg_weight_9_45;
wire signed[31:0]    reg_psum_9_45;
wire signed[31:0]    reg_weight_9_46;
wire signed[31:0]    reg_psum_9_46;
wire signed[31:0]    reg_weight_9_47;
wire signed[31:0]    reg_psum_9_47;
wire signed[31:0]    reg_weight_9_48;
wire signed[31:0]    reg_psum_9_48;
wire signed[31:0]    reg_weight_9_49;
wire signed[31:0]    reg_psum_9_49;
wire signed[31:0]    reg_weight_9_50;
wire signed[31:0]    reg_psum_9_50;
wire signed[31:0]    reg_weight_9_51;
wire signed[31:0]    reg_psum_9_51;
wire signed[31:0]    reg_weight_9_52;
wire signed[31:0]    reg_psum_9_52;
wire signed[31:0]    reg_weight_9_53;
wire signed[31:0]    reg_psum_9_53;
wire signed[31:0]    reg_weight_9_54;
wire signed[31:0]    reg_psum_9_54;
wire signed[31:0]    reg_weight_9_55;
wire signed[31:0]    reg_psum_9_55;
wire signed[31:0]    reg_weight_9_56;
wire signed[31:0]    reg_psum_9_56;
wire signed[31:0]    reg_weight_9_57;
wire signed[31:0]    reg_psum_9_57;
wire signed[31:0]    reg_weight_9_58;
wire signed[31:0]    reg_psum_9_58;
wire signed[31:0]    reg_weight_9_59;
wire signed[31:0]    reg_psum_9_59;
wire signed[31:0]    reg_weight_9_60;
wire signed[31:0]    reg_psum_9_60;
wire signed[31:0]    reg_weight_9_61;
wire signed[31:0]    reg_psum_9_61;
wire signed[31:0]    reg_weight_9_62;
wire signed[31:0]    reg_psum_9_62;
wire signed[31:0]    reg_weight_9_63;
wire signed[31:0]    reg_psum_9_63;
wire signed[31:0]    reg_weight_10_0;
wire signed[31:0]    reg_psum_10_0;
wire signed[31:0]    reg_weight_10_1;
wire signed[31:0]    reg_psum_10_1;
wire signed[31:0]    reg_weight_10_2;
wire signed[31:0]    reg_psum_10_2;
wire signed[31:0]    reg_weight_10_3;
wire signed[31:0]    reg_psum_10_3;
wire signed[31:0]    reg_weight_10_4;
wire signed[31:0]    reg_psum_10_4;
wire signed[31:0]    reg_weight_10_5;
wire signed[31:0]    reg_psum_10_5;
wire signed[31:0]    reg_weight_10_6;
wire signed[31:0]    reg_psum_10_6;
wire signed[31:0]    reg_weight_10_7;
wire signed[31:0]    reg_psum_10_7;
wire signed[31:0]    reg_weight_10_8;
wire signed[31:0]    reg_psum_10_8;
wire signed[31:0]    reg_weight_10_9;
wire signed[31:0]    reg_psum_10_9;
wire signed[31:0]    reg_weight_10_10;
wire signed[31:0]    reg_psum_10_10;
wire signed[31:0]    reg_weight_10_11;
wire signed[31:0]    reg_psum_10_11;
wire signed[31:0]    reg_weight_10_12;
wire signed[31:0]    reg_psum_10_12;
wire signed[31:0]    reg_weight_10_13;
wire signed[31:0]    reg_psum_10_13;
wire signed[31:0]    reg_weight_10_14;
wire signed[31:0]    reg_psum_10_14;
wire signed[31:0]    reg_weight_10_15;
wire signed[31:0]    reg_psum_10_15;
wire signed[31:0]    reg_weight_10_16;
wire signed[31:0]    reg_psum_10_16;
wire signed[31:0]    reg_weight_10_17;
wire signed[31:0]    reg_psum_10_17;
wire signed[31:0]    reg_weight_10_18;
wire signed[31:0]    reg_psum_10_18;
wire signed[31:0]    reg_weight_10_19;
wire signed[31:0]    reg_psum_10_19;
wire signed[31:0]    reg_weight_10_20;
wire signed[31:0]    reg_psum_10_20;
wire signed[31:0]    reg_weight_10_21;
wire signed[31:0]    reg_psum_10_21;
wire signed[31:0]    reg_weight_10_22;
wire signed[31:0]    reg_psum_10_22;
wire signed[31:0]    reg_weight_10_23;
wire signed[31:0]    reg_psum_10_23;
wire signed[31:0]    reg_weight_10_24;
wire signed[31:0]    reg_psum_10_24;
wire signed[31:0]    reg_weight_10_25;
wire signed[31:0]    reg_psum_10_25;
wire signed[31:0]    reg_weight_10_26;
wire signed[31:0]    reg_psum_10_26;
wire signed[31:0]    reg_weight_10_27;
wire signed[31:0]    reg_psum_10_27;
wire signed[31:0]    reg_weight_10_28;
wire signed[31:0]    reg_psum_10_28;
wire signed[31:0]    reg_weight_10_29;
wire signed[31:0]    reg_psum_10_29;
wire signed[31:0]    reg_weight_10_30;
wire signed[31:0]    reg_psum_10_30;
wire signed[31:0]    reg_weight_10_31;
wire signed[31:0]    reg_psum_10_31;
wire signed[31:0]    reg_weight_10_32;
wire signed[31:0]    reg_psum_10_32;
wire signed[31:0]    reg_weight_10_33;
wire signed[31:0]    reg_psum_10_33;
wire signed[31:0]    reg_weight_10_34;
wire signed[31:0]    reg_psum_10_34;
wire signed[31:0]    reg_weight_10_35;
wire signed[31:0]    reg_psum_10_35;
wire signed[31:0]    reg_weight_10_36;
wire signed[31:0]    reg_psum_10_36;
wire signed[31:0]    reg_weight_10_37;
wire signed[31:0]    reg_psum_10_37;
wire signed[31:0]    reg_weight_10_38;
wire signed[31:0]    reg_psum_10_38;
wire signed[31:0]    reg_weight_10_39;
wire signed[31:0]    reg_psum_10_39;
wire signed[31:0]    reg_weight_10_40;
wire signed[31:0]    reg_psum_10_40;
wire signed[31:0]    reg_weight_10_41;
wire signed[31:0]    reg_psum_10_41;
wire signed[31:0]    reg_weight_10_42;
wire signed[31:0]    reg_psum_10_42;
wire signed[31:0]    reg_weight_10_43;
wire signed[31:0]    reg_psum_10_43;
wire signed[31:0]    reg_weight_10_44;
wire signed[31:0]    reg_psum_10_44;
wire signed[31:0]    reg_weight_10_45;
wire signed[31:0]    reg_psum_10_45;
wire signed[31:0]    reg_weight_10_46;
wire signed[31:0]    reg_psum_10_46;
wire signed[31:0]    reg_weight_10_47;
wire signed[31:0]    reg_psum_10_47;
wire signed[31:0]    reg_weight_10_48;
wire signed[31:0]    reg_psum_10_48;
wire signed[31:0]    reg_weight_10_49;
wire signed[31:0]    reg_psum_10_49;
wire signed[31:0]    reg_weight_10_50;
wire signed[31:0]    reg_psum_10_50;
wire signed[31:0]    reg_weight_10_51;
wire signed[31:0]    reg_psum_10_51;
wire signed[31:0]    reg_weight_10_52;
wire signed[31:0]    reg_psum_10_52;
wire signed[31:0]    reg_weight_10_53;
wire signed[31:0]    reg_psum_10_53;
wire signed[31:0]    reg_weight_10_54;
wire signed[31:0]    reg_psum_10_54;
wire signed[31:0]    reg_weight_10_55;
wire signed[31:0]    reg_psum_10_55;
wire signed[31:0]    reg_weight_10_56;
wire signed[31:0]    reg_psum_10_56;
wire signed[31:0]    reg_weight_10_57;
wire signed[31:0]    reg_psum_10_57;
wire signed[31:0]    reg_weight_10_58;
wire signed[31:0]    reg_psum_10_58;
wire signed[31:0]    reg_weight_10_59;
wire signed[31:0]    reg_psum_10_59;
wire signed[31:0]    reg_weight_10_60;
wire signed[31:0]    reg_psum_10_60;
wire signed[31:0]    reg_weight_10_61;
wire signed[31:0]    reg_psum_10_61;
wire signed[31:0]    reg_weight_10_62;
wire signed[31:0]    reg_psum_10_62;
wire signed[31:0]    reg_weight_10_63;
wire signed[31:0]    reg_psum_10_63;
wire signed[31:0]    reg_weight_11_0;
wire signed[31:0]    reg_psum_11_0;
wire signed[31:0]    reg_weight_11_1;
wire signed[31:0]    reg_psum_11_1;
wire signed[31:0]    reg_weight_11_2;
wire signed[31:0]    reg_psum_11_2;
wire signed[31:0]    reg_weight_11_3;
wire signed[31:0]    reg_psum_11_3;
wire signed[31:0]    reg_weight_11_4;
wire signed[31:0]    reg_psum_11_4;
wire signed[31:0]    reg_weight_11_5;
wire signed[31:0]    reg_psum_11_5;
wire signed[31:0]    reg_weight_11_6;
wire signed[31:0]    reg_psum_11_6;
wire signed[31:0]    reg_weight_11_7;
wire signed[31:0]    reg_psum_11_7;
wire signed[31:0]    reg_weight_11_8;
wire signed[31:0]    reg_psum_11_8;
wire signed[31:0]    reg_weight_11_9;
wire signed[31:0]    reg_psum_11_9;
wire signed[31:0]    reg_weight_11_10;
wire signed[31:0]    reg_psum_11_10;
wire signed[31:0]    reg_weight_11_11;
wire signed[31:0]    reg_psum_11_11;
wire signed[31:0]    reg_weight_11_12;
wire signed[31:0]    reg_psum_11_12;
wire signed[31:0]    reg_weight_11_13;
wire signed[31:0]    reg_psum_11_13;
wire signed[31:0]    reg_weight_11_14;
wire signed[31:0]    reg_psum_11_14;
wire signed[31:0]    reg_weight_11_15;
wire signed[31:0]    reg_psum_11_15;
wire signed[31:0]    reg_weight_11_16;
wire signed[31:0]    reg_psum_11_16;
wire signed[31:0]    reg_weight_11_17;
wire signed[31:0]    reg_psum_11_17;
wire signed[31:0]    reg_weight_11_18;
wire signed[31:0]    reg_psum_11_18;
wire signed[31:0]    reg_weight_11_19;
wire signed[31:0]    reg_psum_11_19;
wire signed[31:0]    reg_weight_11_20;
wire signed[31:0]    reg_psum_11_20;
wire signed[31:0]    reg_weight_11_21;
wire signed[31:0]    reg_psum_11_21;
wire signed[31:0]    reg_weight_11_22;
wire signed[31:0]    reg_psum_11_22;
wire signed[31:0]    reg_weight_11_23;
wire signed[31:0]    reg_psum_11_23;
wire signed[31:0]    reg_weight_11_24;
wire signed[31:0]    reg_psum_11_24;
wire signed[31:0]    reg_weight_11_25;
wire signed[31:0]    reg_psum_11_25;
wire signed[31:0]    reg_weight_11_26;
wire signed[31:0]    reg_psum_11_26;
wire signed[31:0]    reg_weight_11_27;
wire signed[31:0]    reg_psum_11_27;
wire signed[31:0]    reg_weight_11_28;
wire signed[31:0]    reg_psum_11_28;
wire signed[31:0]    reg_weight_11_29;
wire signed[31:0]    reg_psum_11_29;
wire signed[31:0]    reg_weight_11_30;
wire signed[31:0]    reg_psum_11_30;
wire signed[31:0]    reg_weight_11_31;
wire signed[31:0]    reg_psum_11_31;
wire signed[31:0]    reg_weight_11_32;
wire signed[31:0]    reg_psum_11_32;
wire signed[31:0]    reg_weight_11_33;
wire signed[31:0]    reg_psum_11_33;
wire signed[31:0]    reg_weight_11_34;
wire signed[31:0]    reg_psum_11_34;
wire signed[31:0]    reg_weight_11_35;
wire signed[31:0]    reg_psum_11_35;
wire signed[31:0]    reg_weight_11_36;
wire signed[31:0]    reg_psum_11_36;
wire signed[31:0]    reg_weight_11_37;
wire signed[31:0]    reg_psum_11_37;
wire signed[31:0]    reg_weight_11_38;
wire signed[31:0]    reg_psum_11_38;
wire signed[31:0]    reg_weight_11_39;
wire signed[31:0]    reg_psum_11_39;
wire signed[31:0]    reg_weight_11_40;
wire signed[31:0]    reg_psum_11_40;
wire signed[31:0]    reg_weight_11_41;
wire signed[31:0]    reg_psum_11_41;
wire signed[31:0]    reg_weight_11_42;
wire signed[31:0]    reg_psum_11_42;
wire signed[31:0]    reg_weight_11_43;
wire signed[31:0]    reg_psum_11_43;
wire signed[31:0]    reg_weight_11_44;
wire signed[31:0]    reg_psum_11_44;
wire signed[31:0]    reg_weight_11_45;
wire signed[31:0]    reg_psum_11_45;
wire signed[31:0]    reg_weight_11_46;
wire signed[31:0]    reg_psum_11_46;
wire signed[31:0]    reg_weight_11_47;
wire signed[31:0]    reg_psum_11_47;
wire signed[31:0]    reg_weight_11_48;
wire signed[31:0]    reg_psum_11_48;
wire signed[31:0]    reg_weight_11_49;
wire signed[31:0]    reg_psum_11_49;
wire signed[31:0]    reg_weight_11_50;
wire signed[31:0]    reg_psum_11_50;
wire signed[31:0]    reg_weight_11_51;
wire signed[31:0]    reg_psum_11_51;
wire signed[31:0]    reg_weight_11_52;
wire signed[31:0]    reg_psum_11_52;
wire signed[31:0]    reg_weight_11_53;
wire signed[31:0]    reg_psum_11_53;
wire signed[31:0]    reg_weight_11_54;
wire signed[31:0]    reg_psum_11_54;
wire signed[31:0]    reg_weight_11_55;
wire signed[31:0]    reg_psum_11_55;
wire signed[31:0]    reg_weight_11_56;
wire signed[31:0]    reg_psum_11_56;
wire signed[31:0]    reg_weight_11_57;
wire signed[31:0]    reg_psum_11_57;
wire signed[31:0]    reg_weight_11_58;
wire signed[31:0]    reg_psum_11_58;
wire signed[31:0]    reg_weight_11_59;
wire signed[31:0]    reg_psum_11_59;
wire signed[31:0]    reg_weight_11_60;
wire signed[31:0]    reg_psum_11_60;
wire signed[31:0]    reg_weight_11_61;
wire signed[31:0]    reg_psum_11_61;
wire signed[31:0]    reg_weight_11_62;
wire signed[31:0]    reg_psum_11_62;
wire signed[31:0]    reg_weight_11_63;
wire signed[31:0]    reg_psum_11_63;
wire signed[31:0]    reg_weight_12_0;
wire signed[31:0]    reg_psum_12_0;
wire signed[31:0]    reg_weight_12_1;
wire signed[31:0]    reg_psum_12_1;
wire signed[31:0]    reg_weight_12_2;
wire signed[31:0]    reg_psum_12_2;
wire signed[31:0]    reg_weight_12_3;
wire signed[31:0]    reg_psum_12_3;
wire signed[31:0]    reg_weight_12_4;
wire signed[31:0]    reg_psum_12_4;
wire signed[31:0]    reg_weight_12_5;
wire signed[31:0]    reg_psum_12_5;
wire signed[31:0]    reg_weight_12_6;
wire signed[31:0]    reg_psum_12_6;
wire signed[31:0]    reg_weight_12_7;
wire signed[31:0]    reg_psum_12_7;
wire signed[31:0]    reg_weight_12_8;
wire signed[31:0]    reg_psum_12_8;
wire signed[31:0]    reg_weight_12_9;
wire signed[31:0]    reg_psum_12_9;
wire signed[31:0]    reg_weight_12_10;
wire signed[31:0]    reg_psum_12_10;
wire signed[31:0]    reg_weight_12_11;
wire signed[31:0]    reg_psum_12_11;
wire signed[31:0]    reg_weight_12_12;
wire signed[31:0]    reg_psum_12_12;
wire signed[31:0]    reg_weight_12_13;
wire signed[31:0]    reg_psum_12_13;
wire signed[31:0]    reg_weight_12_14;
wire signed[31:0]    reg_psum_12_14;
wire signed[31:0]    reg_weight_12_15;
wire signed[31:0]    reg_psum_12_15;
wire signed[31:0]    reg_weight_12_16;
wire signed[31:0]    reg_psum_12_16;
wire signed[31:0]    reg_weight_12_17;
wire signed[31:0]    reg_psum_12_17;
wire signed[31:0]    reg_weight_12_18;
wire signed[31:0]    reg_psum_12_18;
wire signed[31:0]    reg_weight_12_19;
wire signed[31:0]    reg_psum_12_19;
wire signed[31:0]    reg_weight_12_20;
wire signed[31:0]    reg_psum_12_20;
wire signed[31:0]    reg_weight_12_21;
wire signed[31:0]    reg_psum_12_21;
wire signed[31:0]    reg_weight_12_22;
wire signed[31:0]    reg_psum_12_22;
wire signed[31:0]    reg_weight_12_23;
wire signed[31:0]    reg_psum_12_23;
wire signed[31:0]    reg_weight_12_24;
wire signed[31:0]    reg_psum_12_24;
wire signed[31:0]    reg_weight_12_25;
wire signed[31:0]    reg_psum_12_25;
wire signed[31:0]    reg_weight_12_26;
wire signed[31:0]    reg_psum_12_26;
wire signed[31:0]    reg_weight_12_27;
wire signed[31:0]    reg_psum_12_27;
wire signed[31:0]    reg_weight_12_28;
wire signed[31:0]    reg_psum_12_28;
wire signed[31:0]    reg_weight_12_29;
wire signed[31:0]    reg_psum_12_29;
wire signed[31:0]    reg_weight_12_30;
wire signed[31:0]    reg_psum_12_30;
wire signed[31:0]    reg_weight_12_31;
wire signed[31:0]    reg_psum_12_31;
wire signed[31:0]    reg_weight_12_32;
wire signed[31:0]    reg_psum_12_32;
wire signed[31:0]    reg_weight_12_33;
wire signed[31:0]    reg_psum_12_33;
wire signed[31:0]    reg_weight_12_34;
wire signed[31:0]    reg_psum_12_34;
wire signed[31:0]    reg_weight_12_35;
wire signed[31:0]    reg_psum_12_35;
wire signed[31:0]    reg_weight_12_36;
wire signed[31:0]    reg_psum_12_36;
wire signed[31:0]    reg_weight_12_37;
wire signed[31:0]    reg_psum_12_37;
wire signed[31:0]    reg_weight_12_38;
wire signed[31:0]    reg_psum_12_38;
wire signed[31:0]    reg_weight_12_39;
wire signed[31:0]    reg_psum_12_39;
wire signed[31:0]    reg_weight_12_40;
wire signed[31:0]    reg_psum_12_40;
wire signed[31:0]    reg_weight_12_41;
wire signed[31:0]    reg_psum_12_41;
wire signed[31:0]    reg_weight_12_42;
wire signed[31:0]    reg_psum_12_42;
wire signed[31:0]    reg_weight_12_43;
wire signed[31:0]    reg_psum_12_43;
wire signed[31:0]    reg_weight_12_44;
wire signed[31:0]    reg_psum_12_44;
wire signed[31:0]    reg_weight_12_45;
wire signed[31:0]    reg_psum_12_45;
wire signed[31:0]    reg_weight_12_46;
wire signed[31:0]    reg_psum_12_46;
wire signed[31:0]    reg_weight_12_47;
wire signed[31:0]    reg_psum_12_47;
wire signed[31:0]    reg_weight_12_48;
wire signed[31:0]    reg_psum_12_48;
wire signed[31:0]    reg_weight_12_49;
wire signed[31:0]    reg_psum_12_49;
wire signed[31:0]    reg_weight_12_50;
wire signed[31:0]    reg_psum_12_50;
wire signed[31:0]    reg_weight_12_51;
wire signed[31:0]    reg_psum_12_51;
wire signed[31:0]    reg_weight_12_52;
wire signed[31:0]    reg_psum_12_52;
wire signed[31:0]    reg_weight_12_53;
wire signed[31:0]    reg_psum_12_53;
wire signed[31:0]    reg_weight_12_54;
wire signed[31:0]    reg_psum_12_54;
wire signed[31:0]    reg_weight_12_55;
wire signed[31:0]    reg_psum_12_55;
wire signed[31:0]    reg_weight_12_56;
wire signed[31:0]    reg_psum_12_56;
wire signed[31:0]    reg_weight_12_57;
wire signed[31:0]    reg_psum_12_57;
wire signed[31:0]    reg_weight_12_58;
wire signed[31:0]    reg_psum_12_58;
wire signed[31:0]    reg_weight_12_59;
wire signed[31:0]    reg_psum_12_59;
wire signed[31:0]    reg_weight_12_60;
wire signed[31:0]    reg_psum_12_60;
wire signed[31:0]    reg_weight_12_61;
wire signed[31:0]    reg_psum_12_61;
wire signed[31:0]    reg_weight_12_62;
wire signed[31:0]    reg_psum_12_62;
wire signed[31:0]    reg_weight_12_63;
wire signed[31:0]    reg_psum_12_63;
wire signed[31:0]    reg_weight_13_0;
wire signed[31:0]    reg_psum_13_0;
wire signed[31:0]    reg_weight_13_1;
wire signed[31:0]    reg_psum_13_1;
wire signed[31:0]    reg_weight_13_2;
wire signed[31:0]    reg_psum_13_2;
wire signed[31:0]    reg_weight_13_3;
wire signed[31:0]    reg_psum_13_3;
wire signed[31:0]    reg_weight_13_4;
wire signed[31:0]    reg_psum_13_4;
wire signed[31:0]    reg_weight_13_5;
wire signed[31:0]    reg_psum_13_5;
wire signed[31:0]    reg_weight_13_6;
wire signed[31:0]    reg_psum_13_6;
wire signed[31:0]    reg_weight_13_7;
wire signed[31:0]    reg_psum_13_7;
wire signed[31:0]    reg_weight_13_8;
wire signed[31:0]    reg_psum_13_8;
wire signed[31:0]    reg_weight_13_9;
wire signed[31:0]    reg_psum_13_9;
wire signed[31:0]    reg_weight_13_10;
wire signed[31:0]    reg_psum_13_10;
wire signed[31:0]    reg_weight_13_11;
wire signed[31:0]    reg_psum_13_11;
wire signed[31:0]    reg_weight_13_12;
wire signed[31:0]    reg_psum_13_12;
wire signed[31:0]    reg_weight_13_13;
wire signed[31:0]    reg_psum_13_13;
wire signed[31:0]    reg_weight_13_14;
wire signed[31:0]    reg_psum_13_14;
wire signed[31:0]    reg_weight_13_15;
wire signed[31:0]    reg_psum_13_15;
wire signed[31:0]    reg_weight_13_16;
wire signed[31:0]    reg_psum_13_16;
wire signed[31:0]    reg_weight_13_17;
wire signed[31:0]    reg_psum_13_17;
wire signed[31:0]    reg_weight_13_18;
wire signed[31:0]    reg_psum_13_18;
wire signed[31:0]    reg_weight_13_19;
wire signed[31:0]    reg_psum_13_19;
wire signed[31:0]    reg_weight_13_20;
wire signed[31:0]    reg_psum_13_20;
wire signed[31:0]    reg_weight_13_21;
wire signed[31:0]    reg_psum_13_21;
wire signed[31:0]    reg_weight_13_22;
wire signed[31:0]    reg_psum_13_22;
wire signed[31:0]    reg_weight_13_23;
wire signed[31:0]    reg_psum_13_23;
wire signed[31:0]    reg_weight_13_24;
wire signed[31:0]    reg_psum_13_24;
wire signed[31:0]    reg_weight_13_25;
wire signed[31:0]    reg_psum_13_25;
wire signed[31:0]    reg_weight_13_26;
wire signed[31:0]    reg_psum_13_26;
wire signed[31:0]    reg_weight_13_27;
wire signed[31:0]    reg_psum_13_27;
wire signed[31:0]    reg_weight_13_28;
wire signed[31:0]    reg_psum_13_28;
wire signed[31:0]    reg_weight_13_29;
wire signed[31:0]    reg_psum_13_29;
wire signed[31:0]    reg_weight_13_30;
wire signed[31:0]    reg_psum_13_30;
wire signed[31:0]    reg_weight_13_31;
wire signed[31:0]    reg_psum_13_31;
wire signed[31:0]    reg_weight_13_32;
wire signed[31:0]    reg_psum_13_32;
wire signed[31:0]    reg_weight_13_33;
wire signed[31:0]    reg_psum_13_33;
wire signed[31:0]    reg_weight_13_34;
wire signed[31:0]    reg_psum_13_34;
wire signed[31:0]    reg_weight_13_35;
wire signed[31:0]    reg_psum_13_35;
wire signed[31:0]    reg_weight_13_36;
wire signed[31:0]    reg_psum_13_36;
wire signed[31:0]    reg_weight_13_37;
wire signed[31:0]    reg_psum_13_37;
wire signed[31:0]    reg_weight_13_38;
wire signed[31:0]    reg_psum_13_38;
wire signed[31:0]    reg_weight_13_39;
wire signed[31:0]    reg_psum_13_39;
wire signed[31:0]    reg_weight_13_40;
wire signed[31:0]    reg_psum_13_40;
wire signed[31:0]    reg_weight_13_41;
wire signed[31:0]    reg_psum_13_41;
wire signed[31:0]    reg_weight_13_42;
wire signed[31:0]    reg_psum_13_42;
wire signed[31:0]    reg_weight_13_43;
wire signed[31:0]    reg_psum_13_43;
wire signed[31:0]    reg_weight_13_44;
wire signed[31:0]    reg_psum_13_44;
wire signed[31:0]    reg_weight_13_45;
wire signed[31:0]    reg_psum_13_45;
wire signed[31:0]    reg_weight_13_46;
wire signed[31:0]    reg_psum_13_46;
wire signed[31:0]    reg_weight_13_47;
wire signed[31:0]    reg_psum_13_47;
wire signed[31:0]    reg_weight_13_48;
wire signed[31:0]    reg_psum_13_48;
wire signed[31:0]    reg_weight_13_49;
wire signed[31:0]    reg_psum_13_49;
wire signed[31:0]    reg_weight_13_50;
wire signed[31:0]    reg_psum_13_50;
wire signed[31:0]    reg_weight_13_51;
wire signed[31:0]    reg_psum_13_51;
wire signed[31:0]    reg_weight_13_52;
wire signed[31:0]    reg_psum_13_52;
wire signed[31:0]    reg_weight_13_53;
wire signed[31:0]    reg_psum_13_53;
wire signed[31:0]    reg_weight_13_54;
wire signed[31:0]    reg_psum_13_54;
wire signed[31:0]    reg_weight_13_55;
wire signed[31:0]    reg_psum_13_55;
wire signed[31:0]    reg_weight_13_56;
wire signed[31:0]    reg_psum_13_56;
wire signed[31:0]    reg_weight_13_57;
wire signed[31:0]    reg_psum_13_57;
wire signed[31:0]    reg_weight_13_58;
wire signed[31:0]    reg_psum_13_58;
wire signed[31:0]    reg_weight_13_59;
wire signed[31:0]    reg_psum_13_59;
wire signed[31:0]    reg_weight_13_60;
wire signed[31:0]    reg_psum_13_60;
wire signed[31:0]    reg_weight_13_61;
wire signed[31:0]    reg_psum_13_61;
wire signed[31:0]    reg_weight_13_62;
wire signed[31:0]    reg_psum_13_62;
wire signed[31:0]    reg_weight_13_63;
wire signed[31:0]    reg_psum_13_63;
wire signed[31:0]    reg_weight_14_0;
wire signed[31:0]    reg_psum_14_0;
wire signed[31:0]    reg_weight_14_1;
wire signed[31:0]    reg_psum_14_1;
wire signed[31:0]    reg_weight_14_2;
wire signed[31:0]    reg_psum_14_2;
wire signed[31:0]    reg_weight_14_3;
wire signed[31:0]    reg_psum_14_3;
wire signed[31:0]    reg_weight_14_4;
wire signed[31:0]    reg_psum_14_4;
wire signed[31:0]    reg_weight_14_5;
wire signed[31:0]    reg_psum_14_5;
wire signed[31:0]    reg_weight_14_6;
wire signed[31:0]    reg_psum_14_6;
wire signed[31:0]    reg_weight_14_7;
wire signed[31:0]    reg_psum_14_7;
wire signed[31:0]    reg_weight_14_8;
wire signed[31:0]    reg_psum_14_8;
wire signed[31:0]    reg_weight_14_9;
wire signed[31:0]    reg_psum_14_9;
wire signed[31:0]    reg_weight_14_10;
wire signed[31:0]    reg_psum_14_10;
wire signed[31:0]    reg_weight_14_11;
wire signed[31:0]    reg_psum_14_11;
wire signed[31:0]    reg_weight_14_12;
wire signed[31:0]    reg_psum_14_12;
wire signed[31:0]    reg_weight_14_13;
wire signed[31:0]    reg_psum_14_13;
wire signed[31:0]    reg_weight_14_14;
wire signed[31:0]    reg_psum_14_14;
wire signed[31:0]    reg_weight_14_15;
wire signed[31:0]    reg_psum_14_15;
wire signed[31:0]    reg_weight_14_16;
wire signed[31:0]    reg_psum_14_16;
wire signed[31:0]    reg_weight_14_17;
wire signed[31:0]    reg_psum_14_17;
wire signed[31:0]    reg_weight_14_18;
wire signed[31:0]    reg_psum_14_18;
wire signed[31:0]    reg_weight_14_19;
wire signed[31:0]    reg_psum_14_19;
wire signed[31:0]    reg_weight_14_20;
wire signed[31:0]    reg_psum_14_20;
wire signed[31:0]    reg_weight_14_21;
wire signed[31:0]    reg_psum_14_21;
wire signed[31:0]    reg_weight_14_22;
wire signed[31:0]    reg_psum_14_22;
wire signed[31:0]    reg_weight_14_23;
wire signed[31:0]    reg_psum_14_23;
wire signed[31:0]    reg_weight_14_24;
wire signed[31:0]    reg_psum_14_24;
wire signed[31:0]    reg_weight_14_25;
wire signed[31:0]    reg_psum_14_25;
wire signed[31:0]    reg_weight_14_26;
wire signed[31:0]    reg_psum_14_26;
wire signed[31:0]    reg_weight_14_27;
wire signed[31:0]    reg_psum_14_27;
wire signed[31:0]    reg_weight_14_28;
wire signed[31:0]    reg_psum_14_28;
wire signed[31:0]    reg_weight_14_29;
wire signed[31:0]    reg_psum_14_29;
wire signed[31:0]    reg_weight_14_30;
wire signed[31:0]    reg_psum_14_30;
wire signed[31:0]    reg_weight_14_31;
wire signed[31:0]    reg_psum_14_31;
wire signed[31:0]    reg_weight_14_32;
wire signed[31:0]    reg_psum_14_32;
wire signed[31:0]    reg_weight_14_33;
wire signed[31:0]    reg_psum_14_33;
wire signed[31:0]    reg_weight_14_34;
wire signed[31:0]    reg_psum_14_34;
wire signed[31:0]    reg_weight_14_35;
wire signed[31:0]    reg_psum_14_35;
wire signed[31:0]    reg_weight_14_36;
wire signed[31:0]    reg_psum_14_36;
wire signed[31:0]    reg_weight_14_37;
wire signed[31:0]    reg_psum_14_37;
wire signed[31:0]    reg_weight_14_38;
wire signed[31:0]    reg_psum_14_38;
wire signed[31:0]    reg_weight_14_39;
wire signed[31:0]    reg_psum_14_39;
wire signed[31:0]    reg_weight_14_40;
wire signed[31:0]    reg_psum_14_40;
wire signed[31:0]    reg_weight_14_41;
wire signed[31:0]    reg_psum_14_41;
wire signed[31:0]    reg_weight_14_42;
wire signed[31:0]    reg_psum_14_42;
wire signed[31:0]    reg_weight_14_43;
wire signed[31:0]    reg_psum_14_43;
wire signed[31:0]    reg_weight_14_44;
wire signed[31:0]    reg_psum_14_44;
wire signed[31:0]    reg_weight_14_45;
wire signed[31:0]    reg_psum_14_45;
wire signed[31:0]    reg_weight_14_46;
wire signed[31:0]    reg_psum_14_46;
wire signed[31:0]    reg_weight_14_47;
wire signed[31:0]    reg_psum_14_47;
wire signed[31:0]    reg_weight_14_48;
wire signed[31:0]    reg_psum_14_48;
wire signed[31:0]    reg_weight_14_49;
wire signed[31:0]    reg_psum_14_49;
wire signed[31:0]    reg_weight_14_50;
wire signed[31:0]    reg_psum_14_50;
wire signed[31:0]    reg_weight_14_51;
wire signed[31:0]    reg_psum_14_51;
wire signed[31:0]    reg_weight_14_52;
wire signed[31:0]    reg_psum_14_52;
wire signed[31:0]    reg_weight_14_53;
wire signed[31:0]    reg_psum_14_53;
wire signed[31:0]    reg_weight_14_54;
wire signed[31:0]    reg_psum_14_54;
wire signed[31:0]    reg_weight_14_55;
wire signed[31:0]    reg_psum_14_55;
wire signed[31:0]    reg_weight_14_56;
wire signed[31:0]    reg_psum_14_56;
wire signed[31:0]    reg_weight_14_57;
wire signed[31:0]    reg_psum_14_57;
wire signed[31:0]    reg_weight_14_58;
wire signed[31:0]    reg_psum_14_58;
wire signed[31:0]    reg_weight_14_59;
wire signed[31:0]    reg_psum_14_59;
wire signed[31:0]    reg_weight_14_60;
wire signed[31:0]    reg_psum_14_60;
wire signed[31:0]    reg_weight_14_61;
wire signed[31:0]    reg_psum_14_61;
wire signed[31:0]    reg_weight_14_62;
wire signed[31:0]    reg_psum_14_62;
wire signed[31:0]    reg_weight_14_63;
wire signed[31:0]    reg_psum_14_63;
wire signed[31:0]    reg_weight_15_0;
wire signed[31:0]    reg_psum_15_0;
wire signed[31:0]    reg_weight_15_1;
wire signed[31:0]    reg_psum_15_1;
wire signed[31:0]    reg_weight_15_2;
wire signed[31:0]    reg_psum_15_2;
wire signed[31:0]    reg_weight_15_3;
wire signed[31:0]    reg_psum_15_3;
wire signed[31:0]    reg_weight_15_4;
wire signed[31:0]    reg_psum_15_4;
wire signed[31:0]    reg_weight_15_5;
wire signed[31:0]    reg_psum_15_5;
wire signed[31:0]    reg_weight_15_6;
wire signed[31:0]    reg_psum_15_6;
wire signed[31:0]    reg_weight_15_7;
wire signed[31:0]    reg_psum_15_7;
wire signed[31:0]    reg_weight_15_8;
wire signed[31:0]    reg_psum_15_8;
wire signed[31:0]    reg_weight_15_9;
wire signed[31:0]    reg_psum_15_9;
wire signed[31:0]    reg_weight_15_10;
wire signed[31:0]    reg_psum_15_10;
wire signed[31:0]    reg_weight_15_11;
wire signed[31:0]    reg_psum_15_11;
wire signed[31:0]    reg_weight_15_12;
wire signed[31:0]    reg_psum_15_12;
wire signed[31:0]    reg_weight_15_13;
wire signed[31:0]    reg_psum_15_13;
wire signed[31:0]    reg_weight_15_14;
wire signed[31:0]    reg_psum_15_14;
wire signed[31:0]    reg_weight_15_15;
wire signed[31:0]    reg_psum_15_15;
wire signed[31:0]    reg_weight_15_16;
wire signed[31:0]    reg_psum_15_16;
wire signed[31:0]    reg_weight_15_17;
wire signed[31:0]    reg_psum_15_17;
wire signed[31:0]    reg_weight_15_18;
wire signed[31:0]    reg_psum_15_18;
wire signed[31:0]    reg_weight_15_19;
wire signed[31:0]    reg_psum_15_19;
wire signed[31:0]    reg_weight_15_20;
wire signed[31:0]    reg_psum_15_20;
wire signed[31:0]    reg_weight_15_21;
wire signed[31:0]    reg_psum_15_21;
wire signed[31:0]    reg_weight_15_22;
wire signed[31:0]    reg_psum_15_22;
wire signed[31:0]    reg_weight_15_23;
wire signed[31:0]    reg_psum_15_23;
wire signed[31:0]    reg_weight_15_24;
wire signed[31:0]    reg_psum_15_24;
wire signed[31:0]    reg_weight_15_25;
wire signed[31:0]    reg_psum_15_25;
wire signed[31:0]    reg_weight_15_26;
wire signed[31:0]    reg_psum_15_26;
wire signed[31:0]    reg_weight_15_27;
wire signed[31:0]    reg_psum_15_27;
wire signed[31:0]    reg_weight_15_28;
wire signed[31:0]    reg_psum_15_28;
wire signed[31:0]    reg_weight_15_29;
wire signed[31:0]    reg_psum_15_29;
wire signed[31:0]    reg_weight_15_30;
wire signed[31:0]    reg_psum_15_30;
wire signed[31:0]    reg_weight_15_31;
wire signed[31:0]    reg_psum_15_31;
wire signed[31:0]    reg_weight_15_32;
wire signed[31:0]    reg_psum_15_32;
wire signed[31:0]    reg_weight_15_33;
wire signed[31:0]    reg_psum_15_33;
wire signed[31:0]    reg_weight_15_34;
wire signed[31:0]    reg_psum_15_34;
wire signed[31:0]    reg_weight_15_35;
wire signed[31:0]    reg_psum_15_35;
wire signed[31:0]    reg_weight_15_36;
wire signed[31:0]    reg_psum_15_36;
wire signed[31:0]    reg_weight_15_37;
wire signed[31:0]    reg_psum_15_37;
wire signed[31:0]    reg_weight_15_38;
wire signed[31:0]    reg_psum_15_38;
wire signed[31:0]    reg_weight_15_39;
wire signed[31:0]    reg_psum_15_39;
wire signed[31:0]    reg_weight_15_40;
wire signed[31:0]    reg_psum_15_40;
wire signed[31:0]    reg_weight_15_41;
wire signed[31:0]    reg_psum_15_41;
wire signed[31:0]    reg_weight_15_42;
wire signed[31:0]    reg_psum_15_42;
wire signed[31:0]    reg_weight_15_43;
wire signed[31:0]    reg_psum_15_43;
wire signed[31:0]    reg_weight_15_44;
wire signed[31:0]    reg_psum_15_44;
wire signed[31:0]    reg_weight_15_45;
wire signed[31:0]    reg_psum_15_45;
wire signed[31:0]    reg_weight_15_46;
wire signed[31:0]    reg_psum_15_46;
wire signed[31:0]    reg_weight_15_47;
wire signed[31:0]    reg_psum_15_47;
wire signed[31:0]    reg_weight_15_48;
wire signed[31:0]    reg_psum_15_48;
wire signed[31:0]    reg_weight_15_49;
wire signed[31:0]    reg_psum_15_49;
wire signed[31:0]    reg_weight_15_50;
wire signed[31:0]    reg_psum_15_50;
wire signed[31:0]    reg_weight_15_51;
wire signed[31:0]    reg_psum_15_51;
wire signed[31:0]    reg_weight_15_52;
wire signed[31:0]    reg_psum_15_52;
wire signed[31:0]    reg_weight_15_53;
wire signed[31:0]    reg_psum_15_53;
wire signed[31:0]    reg_weight_15_54;
wire signed[31:0]    reg_psum_15_54;
wire signed[31:0]    reg_weight_15_55;
wire signed[31:0]    reg_psum_15_55;
wire signed[31:0]    reg_weight_15_56;
wire signed[31:0]    reg_psum_15_56;
wire signed[31:0]    reg_weight_15_57;
wire signed[31:0]    reg_psum_15_57;
wire signed[31:0]    reg_weight_15_58;
wire signed[31:0]    reg_psum_15_58;
wire signed[31:0]    reg_weight_15_59;
wire signed[31:0]    reg_psum_15_59;
wire signed[31:0]    reg_weight_15_60;
wire signed[31:0]    reg_psum_15_60;
wire signed[31:0]    reg_weight_15_61;
wire signed[31:0]    reg_psum_15_61;
wire signed[31:0]    reg_weight_15_62;
wire signed[31:0]    reg_psum_15_62;
wire signed[31:0]    reg_weight_15_63;
wire signed[31:0]    reg_psum_15_63;
wire signed[31:0]    reg_weight_16_0;
wire signed[31:0]    reg_psum_16_0;
wire signed[31:0]    reg_weight_16_1;
wire signed[31:0]    reg_psum_16_1;
wire signed[31:0]    reg_weight_16_2;
wire signed[31:0]    reg_psum_16_2;
wire signed[31:0]    reg_weight_16_3;
wire signed[31:0]    reg_psum_16_3;
wire signed[31:0]    reg_weight_16_4;
wire signed[31:0]    reg_psum_16_4;
wire signed[31:0]    reg_weight_16_5;
wire signed[31:0]    reg_psum_16_5;
wire signed[31:0]    reg_weight_16_6;
wire signed[31:0]    reg_psum_16_6;
wire signed[31:0]    reg_weight_16_7;
wire signed[31:0]    reg_psum_16_7;
wire signed[31:0]    reg_weight_16_8;
wire signed[31:0]    reg_psum_16_8;
wire signed[31:0]    reg_weight_16_9;
wire signed[31:0]    reg_psum_16_9;
wire signed[31:0]    reg_weight_16_10;
wire signed[31:0]    reg_psum_16_10;
wire signed[31:0]    reg_weight_16_11;
wire signed[31:0]    reg_psum_16_11;
wire signed[31:0]    reg_weight_16_12;
wire signed[31:0]    reg_psum_16_12;
wire signed[31:0]    reg_weight_16_13;
wire signed[31:0]    reg_psum_16_13;
wire signed[31:0]    reg_weight_16_14;
wire signed[31:0]    reg_psum_16_14;
wire signed[31:0]    reg_weight_16_15;
wire signed[31:0]    reg_psum_16_15;
wire signed[31:0]    reg_weight_16_16;
wire signed[31:0]    reg_psum_16_16;
wire signed[31:0]    reg_weight_16_17;
wire signed[31:0]    reg_psum_16_17;
wire signed[31:0]    reg_weight_16_18;
wire signed[31:0]    reg_psum_16_18;
wire signed[31:0]    reg_weight_16_19;
wire signed[31:0]    reg_psum_16_19;
wire signed[31:0]    reg_weight_16_20;
wire signed[31:0]    reg_psum_16_20;
wire signed[31:0]    reg_weight_16_21;
wire signed[31:0]    reg_psum_16_21;
wire signed[31:0]    reg_weight_16_22;
wire signed[31:0]    reg_psum_16_22;
wire signed[31:0]    reg_weight_16_23;
wire signed[31:0]    reg_psum_16_23;
wire signed[31:0]    reg_weight_16_24;
wire signed[31:0]    reg_psum_16_24;
wire signed[31:0]    reg_weight_16_25;
wire signed[31:0]    reg_psum_16_25;
wire signed[31:0]    reg_weight_16_26;
wire signed[31:0]    reg_psum_16_26;
wire signed[31:0]    reg_weight_16_27;
wire signed[31:0]    reg_psum_16_27;
wire signed[31:0]    reg_weight_16_28;
wire signed[31:0]    reg_psum_16_28;
wire signed[31:0]    reg_weight_16_29;
wire signed[31:0]    reg_psum_16_29;
wire signed[31:0]    reg_weight_16_30;
wire signed[31:0]    reg_psum_16_30;
wire signed[31:0]    reg_weight_16_31;
wire signed[31:0]    reg_psum_16_31;
wire signed[31:0]    reg_weight_16_32;
wire signed[31:0]    reg_psum_16_32;
wire signed[31:0]    reg_weight_16_33;
wire signed[31:0]    reg_psum_16_33;
wire signed[31:0]    reg_weight_16_34;
wire signed[31:0]    reg_psum_16_34;
wire signed[31:0]    reg_weight_16_35;
wire signed[31:0]    reg_psum_16_35;
wire signed[31:0]    reg_weight_16_36;
wire signed[31:0]    reg_psum_16_36;
wire signed[31:0]    reg_weight_16_37;
wire signed[31:0]    reg_psum_16_37;
wire signed[31:0]    reg_weight_16_38;
wire signed[31:0]    reg_psum_16_38;
wire signed[31:0]    reg_weight_16_39;
wire signed[31:0]    reg_psum_16_39;
wire signed[31:0]    reg_weight_16_40;
wire signed[31:0]    reg_psum_16_40;
wire signed[31:0]    reg_weight_16_41;
wire signed[31:0]    reg_psum_16_41;
wire signed[31:0]    reg_weight_16_42;
wire signed[31:0]    reg_psum_16_42;
wire signed[31:0]    reg_weight_16_43;
wire signed[31:0]    reg_psum_16_43;
wire signed[31:0]    reg_weight_16_44;
wire signed[31:0]    reg_psum_16_44;
wire signed[31:0]    reg_weight_16_45;
wire signed[31:0]    reg_psum_16_45;
wire signed[31:0]    reg_weight_16_46;
wire signed[31:0]    reg_psum_16_46;
wire signed[31:0]    reg_weight_16_47;
wire signed[31:0]    reg_psum_16_47;
wire signed[31:0]    reg_weight_16_48;
wire signed[31:0]    reg_psum_16_48;
wire signed[31:0]    reg_weight_16_49;
wire signed[31:0]    reg_psum_16_49;
wire signed[31:0]    reg_weight_16_50;
wire signed[31:0]    reg_psum_16_50;
wire signed[31:0]    reg_weight_16_51;
wire signed[31:0]    reg_psum_16_51;
wire signed[31:0]    reg_weight_16_52;
wire signed[31:0]    reg_psum_16_52;
wire signed[31:0]    reg_weight_16_53;
wire signed[31:0]    reg_psum_16_53;
wire signed[31:0]    reg_weight_16_54;
wire signed[31:0]    reg_psum_16_54;
wire signed[31:0]    reg_weight_16_55;
wire signed[31:0]    reg_psum_16_55;
wire signed[31:0]    reg_weight_16_56;
wire signed[31:0]    reg_psum_16_56;
wire signed[31:0]    reg_weight_16_57;
wire signed[31:0]    reg_psum_16_57;
wire signed[31:0]    reg_weight_16_58;
wire signed[31:0]    reg_psum_16_58;
wire signed[31:0]    reg_weight_16_59;
wire signed[31:0]    reg_psum_16_59;
wire signed[31:0]    reg_weight_16_60;
wire signed[31:0]    reg_psum_16_60;
wire signed[31:0]    reg_weight_16_61;
wire signed[31:0]    reg_psum_16_61;
wire signed[31:0]    reg_weight_16_62;
wire signed[31:0]    reg_psum_16_62;
wire signed[31:0]    reg_weight_16_63;
wire signed[31:0]    reg_psum_16_63;
wire signed[31:0]    reg_weight_17_0;
wire signed[31:0]    reg_psum_17_0;
wire signed[31:0]    reg_weight_17_1;
wire signed[31:0]    reg_psum_17_1;
wire signed[31:0]    reg_weight_17_2;
wire signed[31:0]    reg_psum_17_2;
wire signed[31:0]    reg_weight_17_3;
wire signed[31:0]    reg_psum_17_3;
wire signed[31:0]    reg_weight_17_4;
wire signed[31:0]    reg_psum_17_4;
wire signed[31:0]    reg_weight_17_5;
wire signed[31:0]    reg_psum_17_5;
wire signed[31:0]    reg_weight_17_6;
wire signed[31:0]    reg_psum_17_6;
wire signed[31:0]    reg_weight_17_7;
wire signed[31:0]    reg_psum_17_7;
wire signed[31:0]    reg_weight_17_8;
wire signed[31:0]    reg_psum_17_8;
wire signed[31:0]    reg_weight_17_9;
wire signed[31:0]    reg_psum_17_9;
wire signed[31:0]    reg_weight_17_10;
wire signed[31:0]    reg_psum_17_10;
wire signed[31:0]    reg_weight_17_11;
wire signed[31:0]    reg_psum_17_11;
wire signed[31:0]    reg_weight_17_12;
wire signed[31:0]    reg_psum_17_12;
wire signed[31:0]    reg_weight_17_13;
wire signed[31:0]    reg_psum_17_13;
wire signed[31:0]    reg_weight_17_14;
wire signed[31:0]    reg_psum_17_14;
wire signed[31:0]    reg_weight_17_15;
wire signed[31:0]    reg_psum_17_15;
wire signed[31:0]    reg_weight_17_16;
wire signed[31:0]    reg_psum_17_16;
wire signed[31:0]    reg_weight_17_17;
wire signed[31:0]    reg_psum_17_17;
wire signed[31:0]    reg_weight_17_18;
wire signed[31:0]    reg_psum_17_18;
wire signed[31:0]    reg_weight_17_19;
wire signed[31:0]    reg_psum_17_19;
wire signed[31:0]    reg_weight_17_20;
wire signed[31:0]    reg_psum_17_20;
wire signed[31:0]    reg_weight_17_21;
wire signed[31:0]    reg_psum_17_21;
wire signed[31:0]    reg_weight_17_22;
wire signed[31:0]    reg_psum_17_22;
wire signed[31:0]    reg_weight_17_23;
wire signed[31:0]    reg_psum_17_23;
wire signed[31:0]    reg_weight_17_24;
wire signed[31:0]    reg_psum_17_24;
wire signed[31:0]    reg_weight_17_25;
wire signed[31:0]    reg_psum_17_25;
wire signed[31:0]    reg_weight_17_26;
wire signed[31:0]    reg_psum_17_26;
wire signed[31:0]    reg_weight_17_27;
wire signed[31:0]    reg_psum_17_27;
wire signed[31:0]    reg_weight_17_28;
wire signed[31:0]    reg_psum_17_28;
wire signed[31:0]    reg_weight_17_29;
wire signed[31:0]    reg_psum_17_29;
wire signed[31:0]    reg_weight_17_30;
wire signed[31:0]    reg_psum_17_30;
wire signed[31:0]    reg_weight_17_31;
wire signed[31:0]    reg_psum_17_31;
wire signed[31:0]    reg_weight_17_32;
wire signed[31:0]    reg_psum_17_32;
wire signed[31:0]    reg_weight_17_33;
wire signed[31:0]    reg_psum_17_33;
wire signed[31:0]    reg_weight_17_34;
wire signed[31:0]    reg_psum_17_34;
wire signed[31:0]    reg_weight_17_35;
wire signed[31:0]    reg_psum_17_35;
wire signed[31:0]    reg_weight_17_36;
wire signed[31:0]    reg_psum_17_36;
wire signed[31:0]    reg_weight_17_37;
wire signed[31:0]    reg_psum_17_37;
wire signed[31:0]    reg_weight_17_38;
wire signed[31:0]    reg_psum_17_38;
wire signed[31:0]    reg_weight_17_39;
wire signed[31:0]    reg_psum_17_39;
wire signed[31:0]    reg_weight_17_40;
wire signed[31:0]    reg_psum_17_40;
wire signed[31:0]    reg_weight_17_41;
wire signed[31:0]    reg_psum_17_41;
wire signed[31:0]    reg_weight_17_42;
wire signed[31:0]    reg_psum_17_42;
wire signed[31:0]    reg_weight_17_43;
wire signed[31:0]    reg_psum_17_43;
wire signed[31:0]    reg_weight_17_44;
wire signed[31:0]    reg_psum_17_44;
wire signed[31:0]    reg_weight_17_45;
wire signed[31:0]    reg_psum_17_45;
wire signed[31:0]    reg_weight_17_46;
wire signed[31:0]    reg_psum_17_46;
wire signed[31:0]    reg_weight_17_47;
wire signed[31:0]    reg_psum_17_47;
wire signed[31:0]    reg_weight_17_48;
wire signed[31:0]    reg_psum_17_48;
wire signed[31:0]    reg_weight_17_49;
wire signed[31:0]    reg_psum_17_49;
wire signed[31:0]    reg_weight_17_50;
wire signed[31:0]    reg_psum_17_50;
wire signed[31:0]    reg_weight_17_51;
wire signed[31:0]    reg_psum_17_51;
wire signed[31:0]    reg_weight_17_52;
wire signed[31:0]    reg_psum_17_52;
wire signed[31:0]    reg_weight_17_53;
wire signed[31:0]    reg_psum_17_53;
wire signed[31:0]    reg_weight_17_54;
wire signed[31:0]    reg_psum_17_54;
wire signed[31:0]    reg_weight_17_55;
wire signed[31:0]    reg_psum_17_55;
wire signed[31:0]    reg_weight_17_56;
wire signed[31:0]    reg_psum_17_56;
wire signed[31:0]    reg_weight_17_57;
wire signed[31:0]    reg_psum_17_57;
wire signed[31:0]    reg_weight_17_58;
wire signed[31:0]    reg_psum_17_58;
wire signed[31:0]    reg_weight_17_59;
wire signed[31:0]    reg_psum_17_59;
wire signed[31:0]    reg_weight_17_60;
wire signed[31:0]    reg_psum_17_60;
wire signed[31:0]    reg_weight_17_61;
wire signed[31:0]    reg_psum_17_61;
wire signed[31:0]    reg_weight_17_62;
wire signed[31:0]    reg_psum_17_62;
wire signed[31:0]    reg_weight_17_63;
wire signed[31:0]    reg_psum_17_63;
wire signed[31:0]    reg_weight_18_0;
wire signed[31:0]    reg_psum_18_0;
wire signed[31:0]    reg_weight_18_1;
wire signed[31:0]    reg_psum_18_1;
wire signed[31:0]    reg_weight_18_2;
wire signed[31:0]    reg_psum_18_2;
wire signed[31:0]    reg_weight_18_3;
wire signed[31:0]    reg_psum_18_3;
wire signed[31:0]    reg_weight_18_4;
wire signed[31:0]    reg_psum_18_4;
wire signed[31:0]    reg_weight_18_5;
wire signed[31:0]    reg_psum_18_5;
wire signed[31:0]    reg_weight_18_6;
wire signed[31:0]    reg_psum_18_6;
wire signed[31:0]    reg_weight_18_7;
wire signed[31:0]    reg_psum_18_7;
wire signed[31:0]    reg_weight_18_8;
wire signed[31:0]    reg_psum_18_8;
wire signed[31:0]    reg_weight_18_9;
wire signed[31:0]    reg_psum_18_9;
wire signed[31:0]    reg_weight_18_10;
wire signed[31:0]    reg_psum_18_10;
wire signed[31:0]    reg_weight_18_11;
wire signed[31:0]    reg_psum_18_11;
wire signed[31:0]    reg_weight_18_12;
wire signed[31:0]    reg_psum_18_12;
wire signed[31:0]    reg_weight_18_13;
wire signed[31:0]    reg_psum_18_13;
wire signed[31:0]    reg_weight_18_14;
wire signed[31:0]    reg_psum_18_14;
wire signed[31:0]    reg_weight_18_15;
wire signed[31:0]    reg_psum_18_15;
wire signed[31:0]    reg_weight_18_16;
wire signed[31:0]    reg_psum_18_16;
wire signed[31:0]    reg_weight_18_17;
wire signed[31:0]    reg_psum_18_17;
wire signed[31:0]    reg_weight_18_18;
wire signed[31:0]    reg_psum_18_18;
wire signed[31:0]    reg_weight_18_19;
wire signed[31:0]    reg_psum_18_19;
wire signed[31:0]    reg_weight_18_20;
wire signed[31:0]    reg_psum_18_20;
wire signed[31:0]    reg_weight_18_21;
wire signed[31:0]    reg_psum_18_21;
wire signed[31:0]    reg_weight_18_22;
wire signed[31:0]    reg_psum_18_22;
wire signed[31:0]    reg_weight_18_23;
wire signed[31:0]    reg_psum_18_23;
wire signed[31:0]    reg_weight_18_24;
wire signed[31:0]    reg_psum_18_24;
wire signed[31:0]    reg_weight_18_25;
wire signed[31:0]    reg_psum_18_25;
wire signed[31:0]    reg_weight_18_26;
wire signed[31:0]    reg_psum_18_26;
wire signed[31:0]    reg_weight_18_27;
wire signed[31:0]    reg_psum_18_27;
wire signed[31:0]    reg_weight_18_28;
wire signed[31:0]    reg_psum_18_28;
wire signed[31:0]    reg_weight_18_29;
wire signed[31:0]    reg_psum_18_29;
wire signed[31:0]    reg_weight_18_30;
wire signed[31:0]    reg_psum_18_30;
wire signed[31:0]    reg_weight_18_31;
wire signed[31:0]    reg_psum_18_31;
wire signed[31:0]    reg_weight_18_32;
wire signed[31:0]    reg_psum_18_32;
wire signed[31:0]    reg_weight_18_33;
wire signed[31:0]    reg_psum_18_33;
wire signed[31:0]    reg_weight_18_34;
wire signed[31:0]    reg_psum_18_34;
wire signed[31:0]    reg_weight_18_35;
wire signed[31:0]    reg_psum_18_35;
wire signed[31:0]    reg_weight_18_36;
wire signed[31:0]    reg_psum_18_36;
wire signed[31:0]    reg_weight_18_37;
wire signed[31:0]    reg_psum_18_37;
wire signed[31:0]    reg_weight_18_38;
wire signed[31:0]    reg_psum_18_38;
wire signed[31:0]    reg_weight_18_39;
wire signed[31:0]    reg_psum_18_39;
wire signed[31:0]    reg_weight_18_40;
wire signed[31:0]    reg_psum_18_40;
wire signed[31:0]    reg_weight_18_41;
wire signed[31:0]    reg_psum_18_41;
wire signed[31:0]    reg_weight_18_42;
wire signed[31:0]    reg_psum_18_42;
wire signed[31:0]    reg_weight_18_43;
wire signed[31:0]    reg_psum_18_43;
wire signed[31:0]    reg_weight_18_44;
wire signed[31:0]    reg_psum_18_44;
wire signed[31:0]    reg_weight_18_45;
wire signed[31:0]    reg_psum_18_45;
wire signed[31:0]    reg_weight_18_46;
wire signed[31:0]    reg_psum_18_46;
wire signed[31:0]    reg_weight_18_47;
wire signed[31:0]    reg_psum_18_47;
wire signed[31:0]    reg_weight_18_48;
wire signed[31:0]    reg_psum_18_48;
wire signed[31:0]    reg_weight_18_49;
wire signed[31:0]    reg_psum_18_49;
wire signed[31:0]    reg_weight_18_50;
wire signed[31:0]    reg_psum_18_50;
wire signed[31:0]    reg_weight_18_51;
wire signed[31:0]    reg_psum_18_51;
wire signed[31:0]    reg_weight_18_52;
wire signed[31:0]    reg_psum_18_52;
wire signed[31:0]    reg_weight_18_53;
wire signed[31:0]    reg_psum_18_53;
wire signed[31:0]    reg_weight_18_54;
wire signed[31:0]    reg_psum_18_54;
wire signed[31:0]    reg_weight_18_55;
wire signed[31:0]    reg_psum_18_55;
wire signed[31:0]    reg_weight_18_56;
wire signed[31:0]    reg_psum_18_56;
wire signed[31:0]    reg_weight_18_57;
wire signed[31:0]    reg_psum_18_57;
wire signed[31:0]    reg_weight_18_58;
wire signed[31:0]    reg_psum_18_58;
wire signed[31:0]    reg_weight_18_59;
wire signed[31:0]    reg_psum_18_59;
wire signed[31:0]    reg_weight_18_60;
wire signed[31:0]    reg_psum_18_60;
wire signed[31:0]    reg_weight_18_61;
wire signed[31:0]    reg_psum_18_61;
wire signed[31:0]    reg_weight_18_62;
wire signed[31:0]    reg_psum_18_62;
wire signed[31:0]    reg_weight_18_63;
wire signed[31:0]    reg_psum_18_63;
wire signed[31:0]    reg_weight_19_0;
wire signed[31:0]    reg_psum_19_0;
wire signed[31:0]    reg_weight_19_1;
wire signed[31:0]    reg_psum_19_1;
wire signed[31:0]    reg_weight_19_2;
wire signed[31:0]    reg_psum_19_2;
wire signed[31:0]    reg_weight_19_3;
wire signed[31:0]    reg_psum_19_3;
wire signed[31:0]    reg_weight_19_4;
wire signed[31:0]    reg_psum_19_4;
wire signed[31:0]    reg_weight_19_5;
wire signed[31:0]    reg_psum_19_5;
wire signed[31:0]    reg_weight_19_6;
wire signed[31:0]    reg_psum_19_6;
wire signed[31:0]    reg_weight_19_7;
wire signed[31:0]    reg_psum_19_7;
wire signed[31:0]    reg_weight_19_8;
wire signed[31:0]    reg_psum_19_8;
wire signed[31:0]    reg_weight_19_9;
wire signed[31:0]    reg_psum_19_9;
wire signed[31:0]    reg_weight_19_10;
wire signed[31:0]    reg_psum_19_10;
wire signed[31:0]    reg_weight_19_11;
wire signed[31:0]    reg_psum_19_11;
wire signed[31:0]    reg_weight_19_12;
wire signed[31:0]    reg_psum_19_12;
wire signed[31:0]    reg_weight_19_13;
wire signed[31:0]    reg_psum_19_13;
wire signed[31:0]    reg_weight_19_14;
wire signed[31:0]    reg_psum_19_14;
wire signed[31:0]    reg_weight_19_15;
wire signed[31:0]    reg_psum_19_15;
wire signed[31:0]    reg_weight_19_16;
wire signed[31:0]    reg_psum_19_16;
wire signed[31:0]    reg_weight_19_17;
wire signed[31:0]    reg_psum_19_17;
wire signed[31:0]    reg_weight_19_18;
wire signed[31:0]    reg_psum_19_18;
wire signed[31:0]    reg_weight_19_19;
wire signed[31:0]    reg_psum_19_19;
wire signed[31:0]    reg_weight_19_20;
wire signed[31:0]    reg_psum_19_20;
wire signed[31:0]    reg_weight_19_21;
wire signed[31:0]    reg_psum_19_21;
wire signed[31:0]    reg_weight_19_22;
wire signed[31:0]    reg_psum_19_22;
wire signed[31:0]    reg_weight_19_23;
wire signed[31:0]    reg_psum_19_23;
wire signed[31:0]    reg_weight_19_24;
wire signed[31:0]    reg_psum_19_24;
wire signed[31:0]    reg_weight_19_25;
wire signed[31:0]    reg_psum_19_25;
wire signed[31:0]    reg_weight_19_26;
wire signed[31:0]    reg_psum_19_26;
wire signed[31:0]    reg_weight_19_27;
wire signed[31:0]    reg_psum_19_27;
wire signed[31:0]    reg_weight_19_28;
wire signed[31:0]    reg_psum_19_28;
wire signed[31:0]    reg_weight_19_29;
wire signed[31:0]    reg_psum_19_29;
wire signed[31:0]    reg_weight_19_30;
wire signed[31:0]    reg_psum_19_30;
wire signed[31:0]    reg_weight_19_31;
wire signed[31:0]    reg_psum_19_31;
wire signed[31:0]    reg_weight_19_32;
wire signed[31:0]    reg_psum_19_32;
wire signed[31:0]    reg_weight_19_33;
wire signed[31:0]    reg_psum_19_33;
wire signed[31:0]    reg_weight_19_34;
wire signed[31:0]    reg_psum_19_34;
wire signed[31:0]    reg_weight_19_35;
wire signed[31:0]    reg_psum_19_35;
wire signed[31:0]    reg_weight_19_36;
wire signed[31:0]    reg_psum_19_36;
wire signed[31:0]    reg_weight_19_37;
wire signed[31:0]    reg_psum_19_37;
wire signed[31:0]    reg_weight_19_38;
wire signed[31:0]    reg_psum_19_38;
wire signed[31:0]    reg_weight_19_39;
wire signed[31:0]    reg_psum_19_39;
wire signed[31:0]    reg_weight_19_40;
wire signed[31:0]    reg_psum_19_40;
wire signed[31:0]    reg_weight_19_41;
wire signed[31:0]    reg_psum_19_41;
wire signed[31:0]    reg_weight_19_42;
wire signed[31:0]    reg_psum_19_42;
wire signed[31:0]    reg_weight_19_43;
wire signed[31:0]    reg_psum_19_43;
wire signed[31:0]    reg_weight_19_44;
wire signed[31:0]    reg_psum_19_44;
wire signed[31:0]    reg_weight_19_45;
wire signed[31:0]    reg_psum_19_45;
wire signed[31:0]    reg_weight_19_46;
wire signed[31:0]    reg_psum_19_46;
wire signed[31:0]    reg_weight_19_47;
wire signed[31:0]    reg_psum_19_47;
wire signed[31:0]    reg_weight_19_48;
wire signed[31:0]    reg_psum_19_48;
wire signed[31:0]    reg_weight_19_49;
wire signed[31:0]    reg_psum_19_49;
wire signed[31:0]    reg_weight_19_50;
wire signed[31:0]    reg_psum_19_50;
wire signed[31:0]    reg_weight_19_51;
wire signed[31:0]    reg_psum_19_51;
wire signed[31:0]    reg_weight_19_52;
wire signed[31:0]    reg_psum_19_52;
wire signed[31:0]    reg_weight_19_53;
wire signed[31:0]    reg_psum_19_53;
wire signed[31:0]    reg_weight_19_54;
wire signed[31:0]    reg_psum_19_54;
wire signed[31:0]    reg_weight_19_55;
wire signed[31:0]    reg_psum_19_55;
wire signed[31:0]    reg_weight_19_56;
wire signed[31:0]    reg_psum_19_56;
wire signed[31:0]    reg_weight_19_57;
wire signed[31:0]    reg_psum_19_57;
wire signed[31:0]    reg_weight_19_58;
wire signed[31:0]    reg_psum_19_58;
wire signed[31:0]    reg_weight_19_59;
wire signed[31:0]    reg_psum_19_59;
wire signed[31:0]    reg_weight_19_60;
wire signed[31:0]    reg_psum_19_60;
wire signed[31:0]    reg_weight_19_61;
wire signed[31:0]    reg_psum_19_61;
wire signed[31:0]    reg_weight_19_62;
wire signed[31:0]    reg_psum_19_62;
wire signed[31:0]    reg_weight_19_63;
wire signed[31:0]    reg_psum_19_63;
wire signed[31:0]    reg_weight_20_0;
wire signed[31:0]    reg_psum_20_0;
wire signed[31:0]    reg_weight_20_1;
wire signed[31:0]    reg_psum_20_1;
wire signed[31:0]    reg_weight_20_2;
wire signed[31:0]    reg_psum_20_2;
wire signed[31:0]    reg_weight_20_3;
wire signed[31:0]    reg_psum_20_3;
wire signed[31:0]    reg_weight_20_4;
wire signed[31:0]    reg_psum_20_4;
wire signed[31:0]    reg_weight_20_5;
wire signed[31:0]    reg_psum_20_5;
wire signed[31:0]    reg_weight_20_6;
wire signed[31:0]    reg_psum_20_6;
wire signed[31:0]    reg_weight_20_7;
wire signed[31:0]    reg_psum_20_7;
wire signed[31:0]    reg_weight_20_8;
wire signed[31:0]    reg_psum_20_8;
wire signed[31:0]    reg_weight_20_9;
wire signed[31:0]    reg_psum_20_9;
wire signed[31:0]    reg_weight_20_10;
wire signed[31:0]    reg_psum_20_10;
wire signed[31:0]    reg_weight_20_11;
wire signed[31:0]    reg_psum_20_11;
wire signed[31:0]    reg_weight_20_12;
wire signed[31:0]    reg_psum_20_12;
wire signed[31:0]    reg_weight_20_13;
wire signed[31:0]    reg_psum_20_13;
wire signed[31:0]    reg_weight_20_14;
wire signed[31:0]    reg_psum_20_14;
wire signed[31:0]    reg_weight_20_15;
wire signed[31:0]    reg_psum_20_15;
wire signed[31:0]    reg_weight_20_16;
wire signed[31:0]    reg_psum_20_16;
wire signed[31:0]    reg_weight_20_17;
wire signed[31:0]    reg_psum_20_17;
wire signed[31:0]    reg_weight_20_18;
wire signed[31:0]    reg_psum_20_18;
wire signed[31:0]    reg_weight_20_19;
wire signed[31:0]    reg_psum_20_19;
wire signed[31:0]    reg_weight_20_20;
wire signed[31:0]    reg_psum_20_20;
wire signed[31:0]    reg_weight_20_21;
wire signed[31:0]    reg_psum_20_21;
wire signed[31:0]    reg_weight_20_22;
wire signed[31:0]    reg_psum_20_22;
wire signed[31:0]    reg_weight_20_23;
wire signed[31:0]    reg_psum_20_23;
wire signed[31:0]    reg_weight_20_24;
wire signed[31:0]    reg_psum_20_24;
wire signed[31:0]    reg_weight_20_25;
wire signed[31:0]    reg_psum_20_25;
wire signed[31:0]    reg_weight_20_26;
wire signed[31:0]    reg_psum_20_26;
wire signed[31:0]    reg_weight_20_27;
wire signed[31:0]    reg_psum_20_27;
wire signed[31:0]    reg_weight_20_28;
wire signed[31:0]    reg_psum_20_28;
wire signed[31:0]    reg_weight_20_29;
wire signed[31:0]    reg_psum_20_29;
wire signed[31:0]    reg_weight_20_30;
wire signed[31:0]    reg_psum_20_30;
wire signed[31:0]    reg_weight_20_31;
wire signed[31:0]    reg_psum_20_31;
wire signed[31:0]    reg_weight_20_32;
wire signed[31:0]    reg_psum_20_32;
wire signed[31:0]    reg_weight_20_33;
wire signed[31:0]    reg_psum_20_33;
wire signed[31:0]    reg_weight_20_34;
wire signed[31:0]    reg_psum_20_34;
wire signed[31:0]    reg_weight_20_35;
wire signed[31:0]    reg_psum_20_35;
wire signed[31:0]    reg_weight_20_36;
wire signed[31:0]    reg_psum_20_36;
wire signed[31:0]    reg_weight_20_37;
wire signed[31:0]    reg_psum_20_37;
wire signed[31:0]    reg_weight_20_38;
wire signed[31:0]    reg_psum_20_38;
wire signed[31:0]    reg_weight_20_39;
wire signed[31:0]    reg_psum_20_39;
wire signed[31:0]    reg_weight_20_40;
wire signed[31:0]    reg_psum_20_40;
wire signed[31:0]    reg_weight_20_41;
wire signed[31:0]    reg_psum_20_41;
wire signed[31:0]    reg_weight_20_42;
wire signed[31:0]    reg_psum_20_42;
wire signed[31:0]    reg_weight_20_43;
wire signed[31:0]    reg_psum_20_43;
wire signed[31:0]    reg_weight_20_44;
wire signed[31:0]    reg_psum_20_44;
wire signed[31:0]    reg_weight_20_45;
wire signed[31:0]    reg_psum_20_45;
wire signed[31:0]    reg_weight_20_46;
wire signed[31:0]    reg_psum_20_46;
wire signed[31:0]    reg_weight_20_47;
wire signed[31:0]    reg_psum_20_47;
wire signed[31:0]    reg_weight_20_48;
wire signed[31:0]    reg_psum_20_48;
wire signed[31:0]    reg_weight_20_49;
wire signed[31:0]    reg_psum_20_49;
wire signed[31:0]    reg_weight_20_50;
wire signed[31:0]    reg_psum_20_50;
wire signed[31:0]    reg_weight_20_51;
wire signed[31:0]    reg_psum_20_51;
wire signed[31:0]    reg_weight_20_52;
wire signed[31:0]    reg_psum_20_52;
wire signed[31:0]    reg_weight_20_53;
wire signed[31:0]    reg_psum_20_53;
wire signed[31:0]    reg_weight_20_54;
wire signed[31:0]    reg_psum_20_54;
wire signed[31:0]    reg_weight_20_55;
wire signed[31:0]    reg_psum_20_55;
wire signed[31:0]    reg_weight_20_56;
wire signed[31:0]    reg_psum_20_56;
wire signed[31:0]    reg_weight_20_57;
wire signed[31:0]    reg_psum_20_57;
wire signed[31:0]    reg_weight_20_58;
wire signed[31:0]    reg_psum_20_58;
wire signed[31:0]    reg_weight_20_59;
wire signed[31:0]    reg_psum_20_59;
wire signed[31:0]    reg_weight_20_60;
wire signed[31:0]    reg_psum_20_60;
wire signed[31:0]    reg_weight_20_61;
wire signed[31:0]    reg_psum_20_61;
wire signed[31:0]    reg_weight_20_62;
wire signed[31:0]    reg_psum_20_62;
wire signed[31:0]    reg_weight_20_63;
wire signed[31:0]    reg_psum_20_63;
wire signed[31:0]    reg_weight_21_0;
wire signed[31:0]    reg_psum_21_0;
wire signed[31:0]    reg_weight_21_1;
wire signed[31:0]    reg_psum_21_1;
wire signed[31:0]    reg_weight_21_2;
wire signed[31:0]    reg_psum_21_2;
wire signed[31:0]    reg_weight_21_3;
wire signed[31:0]    reg_psum_21_3;
wire signed[31:0]    reg_weight_21_4;
wire signed[31:0]    reg_psum_21_4;
wire signed[31:0]    reg_weight_21_5;
wire signed[31:0]    reg_psum_21_5;
wire signed[31:0]    reg_weight_21_6;
wire signed[31:0]    reg_psum_21_6;
wire signed[31:0]    reg_weight_21_7;
wire signed[31:0]    reg_psum_21_7;
wire signed[31:0]    reg_weight_21_8;
wire signed[31:0]    reg_psum_21_8;
wire signed[31:0]    reg_weight_21_9;
wire signed[31:0]    reg_psum_21_9;
wire signed[31:0]    reg_weight_21_10;
wire signed[31:0]    reg_psum_21_10;
wire signed[31:0]    reg_weight_21_11;
wire signed[31:0]    reg_psum_21_11;
wire signed[31:0]    reg_weight_21_12;
wire signed[31:0]    reg_psum_21_12;
wire signed[31:0]    reg_weight_21_13;
wire signed[31:0]    reg_psum_21_13;
wire signed[31:0]    reg_weight_21_14;
wire signed[31:0]    reg_psum_21_14;
wire signed[31:0]    reg_weight_21_15;
wire signed[31:0]    reg_psum_21_15;
wire signed[31:0]    reg_weight_21_16;
wire signed[31:0]    reg_psum_21_16;
wire signed[31:0]    reg_weight_21_17;
wire signed[31:0]    reg_psum_21_17;
wire signed[31:0]    reg_weight_21_18;
wire signed[31:0]    reg_psum_21_18;
wire signed[31:0]    reg_weight_21_19;
wire signed[31:0]    reg_psum_21_19;
wire signed[31:0]    reg_weight_21_20;
wire signed[31:0]    reg_psum_21_20;
wire signed[31:0]    reg_weight_21_21;
wire signed[31:0]    reg_psum_21_21;
wire signed[31:0]    reg_weight_21_22;
wire signed[31:0]    reg_psum_21_22;
wire signed[31:0]    reg_weight_21_23;
wire signed[31:0]    reg_psum_21_23;
wire signed[31:0]    reg_weight_21_24;
wire signed[31:0]    reg_psum_21_24;
wire signed[31:0]    reg_weight_21_25;
wire signed[31:0]    reg_psum_21_25;
wire signed[31:0]    reg_weight_21_26;
wire signed[31:0]    reg_psum_21_26;
wire signed[31:0]    reg_weight_21_27;
wire signed[31:0]    reg_psum_21_27;
wire signed[31:0]    reg_weight_21_28;
wire signed[31:0]    reg_psum_21_28;
wire signed[31:0]    reg_weight_21_29;
wire signed[31:0]    reg_psum_21_29;
wire signed[31:0]    reg_weight_21_30;
wire signed[31:0]    reg_psum_21_30;
wire signed[31:0]    reg_weight_21_31;
wire signed[31:0]    reg_psum_21_31;
wire signed[31:0]    reg_weight_21_32;
wire signed[31:0]    reg_psum_21_32;
wire signed[31:0]    reg_weight_21_33;
wire signed[31:0]    reg_psum_21_33;
wire signed[31:0]    reg_weight_21_34;
wire signed[31:0]    reg_psum_21_34;
wire signed[31:0]    reg_weight_21_35;
wire signed[31:0]    reg_psum_21_35;
wire signed[31:0]    reg_weight_21_36;
wire signed[31:0]    reg_psum_21_36;
wire signed[31:0]    reg_weight_21_37;
wire signed[31:0]    reg_psum_21_37;
wire signed[31:0]    reg_weight_21_38;
wire signed[31:0]    reg_psum_21_38;
wire signed[31:0]    reg_weight_21_39;
wire signed[31:0]    reg_psum_21_39;
wire signed[31:0]    reg_weight_21_40;
wire signed[31:0]    reg_psum_21_40;
wire signed[31:0]    reg_weight_21_41;
wire signed[31:0]    reg_psum_21_41;
wire signed[31:0]    reg_weight_21_42;
wire signed[31:0]    reg_psum_21_42;
wire signed[31:0]    reg_weight_21_43;
wire signed[31:0]    reg_psum_21_43;
wire signed[31:0]    reg_weight_21_44;
wire signed[31:0]    reg_psum_21_44;
wire signed[31:0]    reg_weight_21_45;
wire signed[31:0]    reg_psum_21_45;
wire signed[31:0]    reg_weight_21_46;
wire signed[31:0]    reg_psum_21_46;
wire signed[31:0]    reg_weight_21_47;
wire signed[31:0]    reg_psum_21_47;
wire signed[31:0]    reg_weight_21_48;
wire signed[31:0]    reg_psum_21_48;
wire signed[31:0]    reg_weight_21_49;
wire signed[31:0]    reg_psum_21_49;
wire signed[31:0]    reg_weight_21_50;
wire signed[31:0]    reg_psum_21_50;
wire signed[31:0]    reg_weight_21_51;
wire signed[31:0]    reg_psum_21_51;
wire signed[31:0]    reg_weight_21_52;
wire signed[31:0]    reg_psum_21_52;
wire signed[31:0]    reg_weight_21_53;
wire signed[31:0]    reg_psum_21_53;
wire signed[31:0]    reg_weight_21_54;
wire signed[31:0]    reg_psum_21_54;
wire signed[31:0]    reg_weight_21_55;
wire signed[31:0]    reg_psum_21_55;
wire signed[31:0]    reg_weight_21_56;
wire signed[31:0]    reg_psum_21_56;
wire signed[31:0]    reg_weight_21_57;
wire signed[31:0]    reg_psum_21_57;
wire signed[31:0]    reg_weight_21_58;
wire signed[31:0]    reg_psum_21_58;
wire signed[31:0]    reg_weight_21_59;
wire signed[31:0]    reg_psum_21_59;
wire signed[31:0]    reg_weight_21_60;
wire signed[31:0]    reg_psum_21_60;
wire signed[31:0]    reg_weight_21_61;
wire signed[31:0]    reg_psum_21_61;
wire signed[31:0]    reg_weight_21_62;
wire signed[31:0]    reg_psum_21_62;
wire signed[31:0]    reg_weight_21_63;
wire signed[31:0]    reg_psum_21_63;
wire signed[31:0]    reg_weight_22_0;
wire signed[31:0]    reg_psum_22_0;
wire signed[31:0]    reg_weight_22_1;
wire signed[31:0]    reg_psum_22_1;
wire signed[31:0]    reg_weight_22_2;
wire signed[31:0]    reg_psum_22_2;
wire signed[31:0]    reg_weight_22_3;
wire signed[31:0]    reg_psum_22_3;
wire signed[31:0]    reg_weight_22_4;
wire signed[31:0]    reg_psum_22_4;
wire signed[31:0]    reg_weight_22_5;
wire signed[31:0]    reg_psum_22_5;
wire signed[31:0]    reg_weight_22_6;
wire signed[31:0]    reg_psum_22_6;
wire signed[31:0]    reg_weight_22_7;
wire signed[31:0]    reg_psum_22_7;
wire signed[31:0]    reg_weight_22_8;
wire signed[31:0]    reg_psum_22_8;
wire signed[31:0]    reg_weight_22_9;
wire signed[31:0]    reg_psum_22_9;
wire signed[31:0]    reg_weight_22_10;
wire signed[31:0]    reg_psum_22_10;
wire signed[31:0]    reg_weight_22_11;
wire signed[31:0]    reg_psum_22_11;
wire signed[31:0]    reg_weight_22_12;
wire signed[31:0]    reg_psum_22_12;
wire signed[31:0]    reg_weight_22_13;
wire signed[31:0]    reg_psum_22_13;
wire signed[31:0]    reg_weight_22_14;
wire signed[31:0]    reg_psum_22_14;
wire signed[31:0]    reg_weight_22_15;
wire signed[31:0]    reg_psum_22_15;
wire signed[31:0]    reg_weight_22_16;
wire signed[31:0]    reg_psum_22_16;
wire signed[31:0]    reg_weight_22_17;
wire signed[31:0]    reg_psum_22_17;
wire signed[31:0]    reg_weight_22_18;
wire signed[31:0]    reg_psum_22_18;
wire signed[31:0]    reg_weight_22_19;
wire signed[31:0]    reg_psum_22_19;
wire signed[31:0]    reg_weight_22_20;
wire signed[31:0]    reg_psum_22_20;
wire signed[31:0]    reg_weight_22_21;
wire signed[31:0]    reg_psum_22_21;
wire signed[31:0]    reg_weight_22_22;
wire signed[31:0]    reg_psum_22_22;
wire signed[31:0]    reg_weight_22_23;
wire signed[31:0]    reg_psum_22_23;
wire signed[31:0]    reg_weight_22_24;
wire signed[31:0]    reg_psum_22_24;
wire signed[31:0]    reg_weight_22_25;
wire signed[31:0]    reg_psum_22_25;
wire signed[31:0]    reg_weight_22_26;
wire signed[31:0]    reg_psum_22_26;
wire signed[31:0]    reg_weight_22_27;
wire signed[31:0]    reg_psum_22_27;
wire signed[31:0]    reg_weight_22_28;
wire signed[31:0]    reg_psum_22_28;
wire signed[31:0]    reg_weight_22_29;
wire signed[31:0]    reg_psum_22_29;
wire signed[31:0]    reg_weight_22_30;
wire signed[31:0]    reg_psum_22_30;
wire signed[31:0]    reg_weight_22_31;
wire signed[31:0]    reg_psum_22_31;
wire signed[31:0]    reg_weight_22_32;
wire signed[31:0]    reg_psum_22_32;
wire signed[31:0]    reg_weight_22_33;
wire signed[31:0]    reg_psum_22_33;
wire signed[31:0]    reg_weight_22_34;
wire signed[31:0]    reg_psum_22_34;
wire signed[31:0]    reg_weight_22_35;
wire signed[31:0]    reg_psum_22_35;
wire signed[31:0]    reg_weight_22_36;
wire signed[31:0]    reg_psum_22_36;
wire signed[31:0]    reg_weight_22_37;
wire signed[31:0]    reg_psum_22_37;
wire signed[31:0]    reg_weight_22_38;
wire signed[31:0]    reg_psum_22_38;
wire signed[31:0]    reg_weight_22_39;
wire signed[31:0]    reg_psum_22_39;
wire signed[31:0]    reg_weight_22_40;
wire signed[31:0]    reg_psum_22_40;
wire signed[31:0]    reg_weight_22_41;
wire signed[31:0]    reg_psum_22_41;
wire signed[31:0]    reg_weight_22_42;
wire signed[31:0]    reg_psum_22_42;
wire signed[31:0]    reg_weight_22_43;
wire signed[31:0]    reg_psum_22_43;
wire signed[31:0]    reg_weight_22_44;
wire signed[31:0]    reg_psum_22_44;
wire signed[31:0]    reg_weight_22_45;
wire signed[31:0]    reg_psum_22_45;
wire signed[31:0]    reg_weight_22_46;
wire signed[31:0]    reg_psum_22_46;
wire signed[31:0]    reg_weight_22_47;
wire signed[31:0]    reg_psum_22_47;
wire signed[31:0]    reg_weight_22_48;
wire signed[31:0]    reg_psum_22_48;
wire signed[31:0]    reg_weight_22_49;
wire signed[31:0]    reg_psum_22_49;
wire signed[31:0]    reg_weight_22_50;
wire signed[31:0]    reg_psum_22_50;
wire signed[31:0]    reg_weight_22_51;
wire signed[31:0]    reg_psum_22_51;
wire signed[31:0]    reg_weight_22_52;
wire signed[31:0]    reg_psum_22_52;
wire signed[31:0]    reg_weight_22_53;
wire signed[31:0]    reg_psum_22_53;
wire signed[31:0]    reg_weight_22_54;
wire signed[31:0]    reg_psum_22_54;
wire signed[31:0]    reg_weight_22_55;
wire signed[31:0]    reg_psum_22_55;
wire signed[31:0]    reg_weight_22_56;
wire signed[31:0]    reg_psum_22_56;
wire signed[31:0]    reg_weight_22_57;
wire signed[31:0]    reg_psum_22_57;
wire signed[31:0]    reg_weight_22_58;
wire signed[31:0]    reg_psum_22_58;
wire signed[31:0]    reg_weight_22_59;
wire signed[31:0]    reg_psum_22_59;
wire signed[31:0]    reg_weight_22_60;
wire signed[31:0]    reg_psum_22_60;
wire signed[31:0]    reg_weight_22_61;
wire signed[31:0]    reg_psum_22_61;
wire signed[31:0]    reg_weight_22_62;
wire signed[31:0]    reg_psum_22_62;
wire signed[31:0]    reg_weight_22_63;
wire signed[31:0]    reg_psum_22_63;
wire signed[31:0]    reg_weight_23_0;
wire signed[31:0]    reg_psum_23_0;
wire signed[31:0]    reg_weight_23_1;
wire signed[31:0]    reg_psum_23_1;
wire signed[31:0]    reg_weight_23_2;
wire signed[31:0]    reg_psum_23_2;
wire signed[31:0]    reg_weight_23_3;
wire signed[31:0]    reg_psum_23_3;
wire signed[31:0]    reg_weight_23_4;
wire signed[31:0]    reg_psum_23_4;
wire signed[31:0]    reg_weight_23_5;
wire signed[31:0]    reg_psum_23_5;
wire signed[31:0]    reg_weight_23_6;
wire signed[31:0]    reg_psum_23_6;
wire signed[31:0]    reg_weight_23_7;
wire signed[31:0]    reg_psum_23_7;
wire signed[31:0]    reg_weight_23_8;
wire signed[31:0]    reg_psum_23_8;
wire signed[31:0]    reg_weight_23_9;
wire signed[31:0]    reg_psum_23_9;
wire signed[31:0]    reg_weight_23_10;
wire signed[31:0]    reg_psum_23_10;
wire signed[31:0]    reg_weight_23_11;
wire signed[31:0]    reg_psum_23_11;
wire signed[31:0]    reg_weight_23_12;
wire signed[31:0]    reg_psum_23_12;
wire signed[31:0]    reg_weight_23_13;
wire signed[31:0]    reg_psum_23_13;
wire signed[31:0]    reg_weight_23_14;
wire signed[31:0]    reg_psum_23_14;
wire signed[31:0]    reg_weight_23_15;
wire signed[31:0]    reg_psum_23_15;
wire signed[31:0]    reg_weight_23_16;
wire signed[31:0]    reg_psum_23_16;
wire signed[31:0]    reg_weight_23_17;
wire signed[31:0]    reg_psum_23_17;
wire signed[31:0]    reg_weight_23_18;
wire signed[31:0]    reg_psum_23_18;
wire signed[31:0]    reg_weight_23_19;
wire signed[31:0]    reg_psum_23_19;
wire signed[31:0]    reg_weight_23_20;
wire signed[31:0]    reg_psum_23_20;
wire signed[31:0]    reg_weight_23_21;
wire signed[31:0]    reg_psum_23_21;
wire signed[31:0]    reg_weight_23_22;
wire signed[31:0]    reg_psum_23_22;
wire signed[31:0]    reg_weight_23_23;
wire signed[31:0]    reg_psum_23_23;
wire signed[31:0]    reg_weight_23_24;
wire signed[31:0]    reg_psum_23_24;
wire signed[31:0]    reg_weight_23_25;
wire signed[31:0]    reg_psum_23_25;
wire signed[31:0]    reg_weight_23_26;
wire signed[31:0]    reg_psum_23_26;
wire signed[31:0]    reg_weight_23_27;
wire signed[31:0]    reg_psum_23_27;
wire signed[31:0]    reg_weight_23_28;
wire signed[31:0]    reg_psum_23_28;
wire signed[31:0]    reg_weight_23_29;
wire signed[31:0]    reg_psum_23_29;
wire signed[31:0]    reg_weight_23_30;
wire signed[31:0]    reg_psum_23_30;
wire signed[31:0]    reg_weight_23_31;
wire signed[31:0]    reg_psum_23_31;
wire signed[31:0]    reg_weight_23_32;
wire signed[31:0]    reg_psum_23_32;
wire signed[31:0]    reg_weight_23_33;
wire signed[31:0]    reg_psum_23_33;
wire signed[31:0]    reg_weight_23_34;
wire signed[31:0]    reg_psum_23_34;
wire signed[31:0]    reg_weight_23_35;
wire signed[31:0]    reg_psum_23_35;
wire signed[31:0]    reg_weight_23_36;
wire signed[31:0]    reg_psum_23_36;
wire signed[31:0]    reg_weight_23_37;
wire signed[31:0]    reg_psum_23_37;
wire signed[31:0]    reg_weight_23_38;
wire signed[31:0]    reg_psum_23_38;
wire signed[31:0]    reg_weight_23_39;
wire signed[31:0]    reg_psum_23_39;
wire signed[31:0]    reg_weight_23_40;
wire signed[31:0]    reg_psum_23_40;
wire signed[31:0]    reg_weight_23_41;
wire signed[31:0]    reg_psum_23_41;
wire signed[31:0]    reg_weight_23_42;
wire signed[31:0]    reg_psum_23_42;
wire signed[31:0]    reg_weight_23_43;
wire signed[31:0]    reg_psum_23_43;
wire signed[31:0]    reg_weight_23_44;
wire signed[31:0]    reg_psum_23_44;
wire signed[31:0]    reg_weight_23_45;
wire signed[31:0]    reg_psum_23_45;
wire signed[31:0]    reg_weight_23_46;
wire signed[31:0]    reg_psum_23_46;
wire signed[31:0]    reg_weight_23_47;
wire signed[31:0]    reg_psum_23_47;
wire signed[31:0]    reg_weight_23_48;
wire signed[31:0]    reg_psum_23_48;
wire signed[31:0]    reg_weight_23_49;
wire signed[31:0]    reg_psum_23_49;
wire signed[31:0]    reg_weight_23_50;
wire signed[31:0]    reg_psum_23_50;
wire signed[31:0]    reg_weight_23_51;
wire signed[31:0]    reg_psum_23_51;
wire signed[31:0]    reg_weight_23_52;
wire signed[31:0]    reg_psum_23_52;
wire signed[31:0]    reg_weight_23_53;
wire signed[31:0]    reg_psum_23_53;
wire signed[31:0]    reg_weight_23_54;
wire signed[31:0]    reg_psum_23_54;
wire signed[31:0]    reg_weight_23_55;
wire signed[31:0]    reg_psum_23_55;
wire signed[31:0]    reg_weight_23_56;
wire signed[31:0]    reg_psum_23_56;
wire signed[31:0]    reg_weight_23_57;
wire signed[31:0]    reg_psum_23_57;
wire signed[31:0]    reg_weight_23_58;
wire signed[31:0]    reg_psum_23_58;
wire signed[31:0]    reg_weight_23_59;
wire signed[31:0]    reg_psum_23_59;
wire signed[31:0]    reg_weight_23_60;
wire signed[31:0]    reg_psum_23_60;
wire signed[31:0]    reg_weight_23_61;
wire signed[31:0]    reg_psum_23_61;
wire signed[31:0]    reg_weight_23_62;
wire signed[31:0]    reg_psum_23_62;
wire signed[31:0]    reg_weight_23_63;
wire signed[31:0]    reg_psum_23_63;
wire signed[31:0]    reg_weight_24_0;
wire signed[31:0]    reg_psum_24_0;
wire signed[31:0]    reg_weight_24_1;
wire signed[31:0]    reg_psum_24_1;
wire signed[31:0]    reg_weight_24_2;
wire signed[31:0]    reg_psum_24_2;
wire signed[31:0]    reg_weight_24_3;
wire signed[31:0]    reg_psum_24_3;
wire signed[31:0]    reg_weight_24_4;
wire signed[31:0]    reg_psum_24_4;
wire signed[31:0]    reg_weight_24_5;
wire signed[31:0]    reg_psum_24_5;
wire signed[31:0]    reg_weight_24_6;
wire signed[31:0]    reg_psum_24_6;
wire signed[31:0]    reg_weight_24_7;
wire signed[31:0]    reg_psum_24_7;
wire signed[31:0]    reg_weight_24_8;
wire signed[31:0]    reg_psum_24_8;
wire signed[31:0]    reg_weight_24_9;
wire signed[31:0]    reg_psum_24_9;
wire signed[31:0]    reg_weight_24_10;
wire signed[31:0]    reg_psum_24_10;
wire signed[31:0]    reg_weight_24_11;
wire signed[31:0]    reg_psum_24_11;
wire signed[31:0]    reg_weight_24_12;
wire signed[31:0]    reg_psum_24_12;
wire signed[31:0]    reg_weight_24_13;
wire signed[31:0]    reg_psum_24_13;
wire signed[31:0]    reg_weight_24_14;
wire signed[31:0]    reg_psum_24_14;
wire signed[31:0]    reg_weight_24_15;
wire signed[31:0]    reg_psum_24_15;
wire signed[31:0]    reg_weight_24_16;
wire signed[31:0]    reg_psum_24_16;
wire signed[31:0]    reg_weight_24_17;
wire signed[31:0]    reg_psum_24_17;
wire signed[31:0]    reg_weight_24_18;
wire signed[31:0]    reg_psum_24_18;
wire signed[31:0]    reg_weight_24_19;
wire signed[31:0]    reg_psum_24_19;
wire signed[31:0]    reg_weight_24_20;
wire signed[31:0]    reg_psum_24_20;
wire signed[31:0]    reg_weight_24_21;
wire signed[31:0]    reg_psum_24_21;
wire signed[31:0]    reg_weight_24_22;
wire signed[31:0]    reg_psum_24_22;
wire signed[31:0]    reg_weight_24_23;
wire signed[31:0]    reg_psum_24_23;
wire signed[31:0]    reg_weight_24_24;
wire signed[31:0]    reg_psum_24_24;
wire signed[31:0]    reg_weight_24_25;
wire signed[31:0]    reg_psum_24_25;
wire signed[31:0]    reg_weight_24_26;
wire signed[31:0]    reg_psum_24_26;
wire signed[31:0]    reg_weight_24_27;
wire signed[31:0]    reg_psum_24_27;
wire signed[31:0]    reg_weight_24_28;
wire signed[31:0]    reg_psum_24_28;
wire signed[31:0]    reg_weight_24_29;
wire signed[31:0]    reg_psum_24_29;
wire signed[31:0]    reg_weight_24_30;
wire signed[31:0]    reg_psum_24_30;
wire signed[31:0]    reg_weight_24_31;
wire signed[31:0]    reg_psum_24_31;
wire signed[31:0]    reg_weight_24_32;
wire signed[31:0]    reg_psum_24_32;
wire signed[31:0]    reg_weight_24_33;
wire signed[31:0]    reg_psum_24_33;
wire signed[31:0]    reg_weight_24_34;
wire signed[31:0]    reg_psum_24_34;
wire signed[31:0]    reg_weight_24_35;
wire signed[31:0]    reg_psum_24_35;
wire signed[31:0]    reg_weight_24_36;
wire signed[31:0]    reg_psum_24_36;
wire signed[31:0]    reg_weight_24_37;
wire signed[31:0]    reg_psum_24_37;
wire signed[31:0]    reg_weight_24_38;
wire signed[31:0]    reg_psum_24_38;
wire signed[31:0]    reg_weight_24_39;
wire signed[31:0]    reg_psum_24_39;
wire signed[31:0]    reg_weight_24_40;
wire signed[31:0]    reg_psum_24_40;
wire signed[31:0]    reg_weight_24_41;
wire signed[31:0]    reg_psum_24_41;
wire signed[31:0]    reg_weight_24_42;
wire signed[31:0]    reg_psum_24_42;
wire signed[31:0]    reg_weight_24_43;
wire signed[31:0]    reg_psum_24_43;
wire signed[31:0]    reg_weight_24_44;
wire signed[31:0]    reg_psum_24_44;
wire signed[31:0]    reg_weight_24_45;
wire signed[31:0]    reg_psum_24_45;
wire signed[31:0]    reg_weight_24_46;
wire signed[31:0]    reg_psum_24_46;
wire signed[31:0]    reg_weight_24_47;
wire signed[31:0]    reg_psum_24_47;
wire signed[31:0]    reg_weight_24_48;
wire signed[31:0]    reg_psum_24_48;
wire signed[31:0]    reg_weight_24_49;
wire signed[31:0]    reg_psum_24_49;
wire signed[31:0]    reg_weight_24_50;
wire signed[31:0]    reg_psum_24_50;
wire signed[31:0]    reg_weight_24_51;
wire signed[31:0]    reg_psum_24_51;
wire signed[31:0]    reg_weight_24_52;
wire signed[31:0]    reg_psum_24_52;
wire signed[31:0]    reg_weight_24_53;
wire signed[31:0]    reg_psum_24_53;
wire signed[31:0]    reg_weight_24_54;
wire signed[31:0]    reg_psum_24_54;
wire signed[31:0]    reg_weight_24_55;
wire signed[31:0]    reg_psum_24_55;
wire signed[31:0]    reg_weight_24_56;
wire signed[31:0]    reg_psum_24_56;
wire signed[31:0]    reg_weight_24_57;
wire signed[31:0]    reg_psum_24_57;
wire signed[31:0]    reg_weight_24_58;
wire signed[31:0]    reg_psum_24_58;
wire signed[31:0]    reg_weight_24_59;
wire signed[31:0]    reg_psum_24_59;
wire signed[31:0]    reg_weight_24_60;
wire signed[31:0]    reg_psum_24_60;
wire signed[31:0]    reg_weight_24_61;
wire signed[31:0]    reg_psum_24_61;
wire signed[31:0]    reg_weight_24_62;
wire signed[31:0]    reg_psum_24_62;
wire signed[31:0]    reg_weight_24_63;
wire signed[31:0]    reg_psum_24_63;
wire signed[31:0]    reg_weight_25_0;
wire signed[31:0]    reg_psum_25_0;
wire signed[31:0]    reg_weight_25_1;
wire signed[31:0]    reg_psum_25_1;
wire signed[31:0]    reg_weight_25_2;
wire signed[31:0]    reg_psum_25_2;
wire signed[31:0]    reg_weight_25_3;
wire signed[31:0]    reg_psum_25_3;
wire signed[31:0]    reg_weight_25_4;
wire signed[31:0]    reg_psum_25_4;
wire signed[31:0]    reg_weight_25_5;
wire signed[31:0]    reg_psum_25_5;
wire signed[31:0]    reg_weight_25_6;
wire signed[31:0]    reg_psum_25_6;
wire signed[31:0]    reg_weight_25_7;
wire signed[31:0]    reg_psum_25_7;
wire signed[31:0]    reg_weight_25_8;
wire signed[31:0]    reg_psum_25_8;
wire signed[31:0]    reg_weight_25_9;
wire signed[31:0]    reg_psum_25_9;
wire signed[31:0]    reg_weight_25_10;
wire signed[31:0]    reg_psum_25_10;
wire signed[31:0]    reg_weight_25_11;
wire signed[31:0]    reg_psum_25_11;
wire signed[31:0]    reg_weight_25_12;
wire signed[31:0]    reg_psum_25_12;
wire signed[31:0]    reg_weight_25_13;
wire signed[31:0]    reg_psum_25_13;
wire signed[31:0]    reg_weight_25_14;
wire signed[31:0]    reg_psum_25_14;
wire signed[31:0]    reg_weight_25_15;
wire signed[31:0]    reg_psum_25_15;
wire signed[31:0]    reg_weight_25_16;
wire signed[31:0]    reg_psum_25_16;
wire signed[31:0]    reg_weight_25_17;
wire signed[31:0]    reg_psum_25_17;
wire signed[31:0]    reg_weight_25_18;
wire signed[31:0]    reg_psum_25_18;
wire signed[31:0]    reg_weight_25_19;
wire signed[31:0]    reg_psum_25_19;
wire signed[31:0]    reg_weight_25_20;
wire signed[31:0]    reg_psum_25_20;
wire signed[31:0]    reg_weight_25_21;
wire signed[31:0]    reg_psum_25_21;
wire signed[31:0]    reg_weight_25_22;
wire signed[31:0]    reg_psum_25_22;
wire signed[31:0]    reg_weight_25_23;
wire signed[31:0]    reg_psum_25_23;
wire signed[31:0]    reg_weight_25_24;
wire signed[31:0]    reg_psum_25_24;
wire signed[31:0]    reg_weight_25_25;
wire signed[31:0]    reg_psum_25_25;
wire signed[31:0]    reg_weight_25_26;
wire signed[31:0]    reg_psum_25_26;
wire signed[31:0]    reg_weight_25_27;
wire signed[31:0]    reg_psum_25_27;
wire signed[31:0]    reg_weight_25_28;
wire signed[31:0]    reg_psum_25_28;
wire signed[31:0]    reg_weight_25_29;
wire signed[31:0]    reg_psum_25_29;
wire signed[31:0]    reg_weight_25_30;
wire signed[31:0]    reg_psum_25_30;
wire signed[31:0]    reg_weight_25_31;
wire signed[31:0]    reg_psum_25_31;
wire signed[31:0]    reg_weight_25_32;
wire signed[31:0]    reg_psum_25_32;
wire signed[31:0]    reg_weight_25_33;
wire signed[31:0]    reg_psum_25_33;
wire signed[31:0]    reg_weight_25_34;
wire signed[31:0]    reg_psum_25_34;
wire signed[31:0]    reg_weight_25_35;
wire signed[31:0]    reg_psum_25_35;
wire signed[31:0]    reg_weight_25_36;
wire signed[31:0]    reg_psum_25_36;
wire signed[31:0]    reg_weight_25_37;
wire signed[31:0]    reg_psum_25_37;
wire signed[31:0]    reg_weight_25_38;
wire signed[31:0]    reg_psum_25_38;
wire signed[31:0]    reg_weight_25_39;
wire signed[31:0]    reg_psum_25_39;
wire signed[31:0]    reg_weight_25_40;
wire signed[31:0]    reg_psum_25_40;
wire signed[31:0]    reg_weight_25_41;
wire signed[31:0]    reg_psum_25_41;
wire signed[31:0]    reg_weight_25_42;
wire signed[31:0]    reg_psum_25_42;
wire signed[31:0]    reg_weight_25_43;
wire signed[31:0]    reg_psum_25_43;
wire signed[31:0]    reg_weight_25_44;
wire signed[31:0]    reg_psum_25_44;
wire signed[31:0]    reg_weight_25_45;
wire signed[31:0]    reg_psum_25_45;
wire signed[31:0]    reg_weight_25_46;
wire signed[31:0]    reg_psum_25_46;
wire signed[31:0]    reg_weight_25_47;
wire signed[31:0]    reg_psum_25_47;
wire signed[31:0]    reg_weight_25_48;
wire signed[31:0]    reg_psum_25_48;
wire signed[31:0]    reg_weight_25_49;
wire signed[31:0]    reg_psum_25_49;
wire signed[31:0]    reg_weight_25_50;
wire signed[31:0]    reg_psum_25_50;
wire signed[31:0]    reg_weight_25_51;
wire signed[31:0]    reg_psum_25_51;
wire signed[31:0]    reg_weight_25_52;
wire signed[31:0]    reg_psum_25_52;
wire signed[31:0]    reg_weight_25_53;
wire signed[31:0]    reg_psum_25_53;
wire signed[31:0]    reg_weight_25_54;
wire signed[31:0]    reg_psum_25_54;
wire signed[31:0]    reg_weight_25_55;
wire signed[31:0]    reg_psum_25_55;
wire signed[31:0]    reg_weight_25_56;
wire signed[31:0]    reg_psum_25_56;
wire signed[31:0]    reg_weight_25_57;
wire signed[31:0]    reg_psum_25_57;
wire signed[31:0]    reg_weight_25_58;
wire signed[31:0]    reg_psum_25_58;
wire signed[31:0]    reg_weight_25_59;
wire signed[31:0]    reg_psum_25_59;
wire signed[31:0]    reg_weight_25_60;
wire signed[31:0]    reg_psum_25_60;
wire signed[31:0]    reg_weight_25_61;
wire signed[31:0]    reg_psum_25_61;
wire signed[31:0]    reg_weight_25_62;
wire signed[31:0]    reg_psum_25_62;
wire signed[31:0]    reg_weight_25_63;
wire signed[31:0]    reg_psum_25_63;
wire signed[31:0]    reg_weight_26_0;
wire signed[31:0]    reg_psum_26_0;
wire signed[31:0]    reg_weight_26_1;
wire signed[31:0]    reg_psum_26_1;
wire signed[31:0]    reg_weight_26_2;
wire signed[31:0]    reg_psum_26_2;
wire signed[31:0]    reg_weight_26_3;
wire signed[31:0]    reg_psum_26_3;
wire signed[31:0]    reg_weight_26_4;
wire signed[31:0]    reg_psum_26_4;
wire signed[31:0]    reg_weight_26_5;
wire signed[31:0]    reg_psum_26_5;
wire signed[31:0]    reg_weight_26_6;
wire signed[31:0]    reg_psum_26_6;
wire signed[31:0]    reg_weight_26_7;
wire signed[31:0]    reg_psum_26_7;
wire signed[31:0]    reg_weight_26_8;
wire signed[31:0]    reg_psum_26_8;
wire signed[31:0]    reg_weight_26_9;
wire signed[31:0]    reg_psum_26_9;
wire signed[31:0]    reg_weight_26_10;
wire signed[31:0]    reg_psum_26_10;
wire signed[31:0]    reg_weight_26_11;
wire signed[31:0]    reg_psum_26_11;
wire signed[31:0]    reg_weight_26_12;
wire signed[31:0]    reg_psum_26_12;
wire signed[31:0]    reg_weight_26_13;
wire signed[31:0]    reg_psum_26_13;
wire signed[31:0]    reg_weight_26_14;
wire signed[31:0]    reg_psum_26_14;
wire signed[31:0]    reg_weight_26_15;
wire signed[31:0]    reg_psum_26_15;
wire signed[31:0]    reg_weight_26_16;
wire signed[31:0]    reg_psum_26_16;
wire signed[31:0]    reg_weight_26_17;
wire signed[31:0]    reg_psum_26_17;
wire signed[31:0]    reg_weight_26_18;
wire signed[31:0]    reg_psum_26_18;
wire signed[31:0]    reg_weight_26_19;
wire signed[31:0]    reg_psum_26_19;
wire signed[31:0]    reg_weight_26_20;
wire signed[31:0]    reg_psum_26_20;
wire signed[31:0]    reg_weight_26_21;
wire signed[31:0]    reg_psum_26_21;
wire signed[31:0]    reg_weight_26_22;
wire signed[31:0]    reg_psum_26_22;
wire signed[31:0]    reg_weight_26_23;
wire signed[31:0]    reg_psum_26_23;
wire signed[31:0]    reg_weight_26_24;
wire signed[31:0]    reg_psum_26_24;
wire signed[31:0]    reg_weight_26_25;
wire signed[31:0]    reg_psum_26_25;
wire signed[31:0]    reg_weight_26_26;
wire signed[31:0]    reg_psum_26_26;
wire signed[31:0]    reg_weight_26_27;
wire signed[31:0]    reg_psum_26_27;
wire signed[31:0]    reg_weight_26_28;
wire signed[31:0]    reg_psum_26_28;
wire signed[31:0]    reg_weight_26_29;
wire signed[31:0]    reg_psum_26_29;
wire signed[31:0]    reg_weight_26_30;
wire signed[31:0]    reg_psum_26_30;
wire signed[31:0]    reg_weight_26_31;
wire signed[31:0]    reg_psum_26_31;
wire signed[31:0]    reg_weight_26_32;
wire signed[31:0]    reg_psum_26_32;
wire signed[31:0]    reg_weight_26_33;
wire signed[31:0]    reg_psum_26_33;
wire signed[31:0]    reg_weight_26_34;
wire signed[31:0]    reg_psum_26_34;
wire signed[31:0]    reg_weight_26_35;
wire signed[31:0]    reg_psum_26_35;
wire signed[31:0]    reg_weight_26_36;
wire signed[31:0]    reg_psum_26_36;
wire signed[31:0]    reg_weight_26_37;
wire signed[31:0]    reg_psum_26_37;
wire signed[31:0]    reg_weight_26_38;
wire signed[31:0]    reg_psum_26_38;
wire signed[31:0]    reg_weight_26_39;
wire signed[31:0]    reg_psum_26_39;
wire signed[31:0]    reg_weight_26_40;
wire signed[31:0]    reg_psum_26_40;
wire signed[31:0]    reg_weight_26_41;
wire signed[31:0]    reg_psum_26_41;
wire signed[31:0]    reg_weight_26_42;
wire signed[31:0]    reg_psum_26_42;
wire signed[31:0]    reg_weight_26_43;
wire signed[31:0]    reg_psum_26_43;
wire signed[31:0]    reg_weight_26_44;
wire signed[31:0]    reg_psum_26_44;
wire signed[31:0]    reg_weight_26_45;
wire signed[31:0]    reg_psum_26_45;
wire signed[31:0]    reg_weight_26_46;
wire signed[31:0]    reg_psum_26_46;
wire signed[31:0]    reg_weight_26_47;
wire signed[31:0]    reg_psum_26_47;
wire signed[31:0]    reg_weight_26_48;
wire signed[31:0]    reg_psum_26_48;
wire signed[31:0]    reg_weight_26_49;
wire signed[31:0]    reg_psum_26_49;
wire signed[31:0]    reg_weight_26_50;
wire signed[31:0]    reg_psum_26_50;
wire signed[31:0]    reg_weight_26_51;
wire signed[31:0]    reg_psum_26_51;
wire signed[31:0]    reg_weight_26_52;
wire signed[31:0]    reg_psum_26_52;
wire signed[31:0]    reg_weight_26_53;
wire signed[31:0]    reg_psum_26_53;
wire signed[31:0]    reg_weight_26_54;
wire signed[31:0]    reg_psum_26_54;
wire signed[31:0]    reg_weight_26_55;
wire signed[31:0]    reg_psum_26_55;
wire signed[31:0]    reg_weight_26_56;
wire signed[31:0]    reg_psum_26_56;
wire signed[31:0]    reg_weight_26_57;
wire signed[31:0]    reg_psum_26_57;
wire signed[31:0]    reg_weight_26_58;
wire signed[31:0]    reg_psum_26_58;
wire signed[31:0]    reg_weight_26_59;
wire signed[31:0]    reg_psum_26_59;
wire signed[31:0]    reg_weight_26_60;
wire signed[31:0]    reg_psum_26_60;
wire signed[31:0]    reg_weight_26_61;
wire signed[31:0]    reg_psum_26_61;
wire signed[31:0]    reg_weight_26_62;
wire signed[31:0]    reg_psum_26_62;
wire signed[31:0]    reg_weight_26_63;
wire signed[31:0]    reg_psum_26_63;
wire signed[31:0]    reg_weight_27_0;
wire signed[31:0]    reg_psum_27_0;
wire signed[31:0]    reg_weight_27_1;
wire signed[31:0]    reg_psum_27_1;
wire signed[31:0]    reg_weight_27_2;
wire signed[31:0]    reg_psum_27_2;
wire signed[31:0]    reg_weight_27_3;
wire signed[31:0]    reg_psum_27_3;
wire signed[31:0]    reg_weight_27_4;
wire signed[31:0]    reg_psum_27_4;
wire signed[31:0]    reg_weight_27_5;
wire signed[31:0]    reg_psum_27_5;
wire signed[31:0]    reg_weight_27_6;
wire signed[31:0]    reg_psum_27_6;
wire signed[31:0]    reg_weight_27_7;
wire signed[31:0]    reg_psum_27_7;
wire signed[31:0]    reg_weight_27_8;
wire signed[31:0]    reg_psum_27_8;
wire signed[31:0]    reg_weight_27_9;
wire signed[31:0]    reg_psum_27_9;
wire signed[31:0]    reg_weight_27_10;
wire signed[31:0]    reg_psum_27_10;
wire signed[31:0]    reg_weight_27_11;
wire signed[31:0]    reg_psum_27_11;
wire signed[31:0]    reg_weight_27_12;
wire signed[31:0]    reg_psum_27_12;
wire signed[31:0]    reg_weight_27_13;
wire signed[31:0]    reg_psum_27_13;
wire signed[31:0]    reg_weight_27_14;
wire signed[31:0]    reg_psum_27_14;
wire signed[31:0]    reg_weight_27_15;
wire signed[31:0]    reg_psum_27_15;
wire signed[31:0]    reg_weight_27_16;
wire signed[31:0]    reg_psum_27_16;
wire signed[31:0]    reg_weight_27_17;
wire signed[31:0]    reg_psum_27_17;
wire signed[31:0]    reg_weight_27_18;
wire signed[31:0]    reg_psum_27_18;
wire signed[31:0]    reg_weight_27_19;
wire signed[31:0]    reg_psum_27_19;
wire signed[31:0]    reg_weight_27_20;
wire signed[31:0]    reg_psum_27_20;
wire signed[31:0]    reg_weight_27_21;
wire signed[31:0]    reg_psum_27_21;
wire signed[31:0]    reg_weight_27_22;
wire signed[31:0]    reg_psum_27_22;
wire signed[31:0]    reg_weight_27_23;
wire signed[31:0]    reg_psum_27_23;
wire signed[31:0]    reg_weight_27_24;
wire signed[31:0]    reg_psum_27_24;
wire signed[31:0]    reg_weight_27_25;
wire signed[31:0]    reg_psum_27_25;
wire signed[31:0]    reg_weight_27_26;
wire signed[31:0]    reg_psum_27_26;
wire signed[31:0]    reg_weight_27_27;
wire signed[31:0]    reg_psum_27_27;
wire signed[31:0]    reg_weight_27_28;
wire signed[31:0]    reg_psum_27_28;
wire signed[31:0]    reg_weight_27_29;
wire signed[31:0]    reg_psum_27_29;
wire signed[31:0]    reg_weight_27_30;
wire signed[31:0]    reg_psum_27_30;
wire signed[31:0]    reg_weight_27_31;
wire signed[31:0]    reg_psum_27_31;
wire signed[31:0]    reg_weight_27_32;
wire signed[31:0]    reg_psum_27_32;
wire signed[31:0]    reg_weight_27_33;
wire signed[31:0]    reg_psum_27_33;
wire signed[31:0]    reg_weight_27_34;
wire signed[31:0]    reg_psum_27_34;
wire signed[31:0]    reg_weight_27_35;
wire signed[31:0]    reg_psum_27_35;
wire signed[31:0]    reg_weight_27_36;
wire signed[31:0]    reg_psum_27_36;
wire signed[31:0]    reg_weight_27_37;
wire signed[31:0]    reg_psum_27_37;
wire signed[31:0]    reg_weight_27_38;
wire signed[31:0]    reg_psum_27_38;
wire signed[31:0]    reg_weight_27_39;
wire signed[31:0]    reg_psum_27_39;
wire signed[31:0]    reg_weight_27_40;
wire signed[31:0]    reg_psum_27_40;
wire signed[31:0]    reg_weight_27_41;
wire signed[31:0]    reg_psum_27_41;
wire signed[31:0]    reg_weight_27_42;
wire signed[31:0]    reg_psum_27_42;
wire signed[31:0]    reg_weight_27_43;
wire signed[31:0]    reg_psum_27_43;
wire signed[31:0]    reg_weight_27_44;
wire signed[31:0]    reg_psum_27_44;
wire signed[31:0]    reg_weight_27_45;
wire signed[31:0]    reg_psum_27_45;
wire signed[31:0]    reg_weight_27_46;
wire signed[31:0]    reg_psum_27_46;
wire signed[31:0]    reg_weight_27_47;
wire signed[31:0]    reg_psum_27_47;
wire signed[31:0]    reg_weight_27_48;
wire signed[31:0]    reg_psum_27_48;
wire signed[31:0]    reg_weight_27_49;
wire signed[31:0]    reg_psum_27_49;
wire signed[31:0]    reg_weight_27_50;
wire signed[31:0]    reg_psum_27_50;
wire signed[31:0]    reg_weight_27_51;
wire signed[31:0]    reg_psum_27_51;
wire signed[31:0]    reg_weight_27_52;
wire signed[31:0]    reg_psum_27_52;
wire signed[31:0]    reg_weight_27_53;
wire signed[31:0]    reg_psum_27_53;
wire signed[31:0]    reg_weight_27_54;
wire signed[31:0]    reg_psum_27_54;
wire signed[31:0]    reg_weight_27_55;
wire signed[31:0]    reg_psum_27_55;
wire signed[31:0]    reg_weight_27_56;
wire signed[31:0]    reg_psum_27_56;
wire signed[31:0]    reg_weight_27_57;
wire signed[31:0]    reg_psum_27_57;
wire signed[31:0]    reg_weight_27_58;
wire signed[31:0]    reg_psum_27_58;
wire signed[31:0]    reg_weight_27_59;
wire signed[31:0]    reg_psum_27_59;
wire signed[31:0]    reg_weight_27_60;
wire signed[31:0]    reg_psum_27_60;
wire signed[31:0]    reg_weight_27_61;
wire signed[31:0]    reg_psum_27_61;
wire signed[31:0]    reg_weight_27_62;
wire signed[31:0]    reg_psum_27_62;
wire signed[31:0]    reg_weight_27_63;
wire signed[31:0]    reg_psum_27_63;
wire signed[31:0]    reg_weight_28_0;
wire signed[31:0]    reg_psum_28_0;
wire signed[31:0]    reg_weight_28_1;
wire signed[31:0]    reg_psum_28_1;
wire signed[31:0]    reg_weight_28_2;
wire signed[31:0]    reg_psum_28_2;
wire signed[31:0]    reg_weight_28_3;
wire signed[31:0]    reg_psum_28_3;
wire signed[31:0]    reg_weight_28_4;
wire signed[31:0]    reg_psum_28_4;
wire signed[31:0]    reg_weight_28_5;
wire signed[31:0]    reg_psum_28_5;
wire signed[31:0]    reg_weight_28_6;
wire signed[31:0]    reg_psum_28_6;
wire signed[31:0]    reg_weight_28_7;
wire signed[31:0]    reg_psum_28_7;
wire signed[31:0]    reg_weight_28_8;
wire signed[31:0]    reg_psum_28_8;
wire signed[31:0]    reg_weight_28_9;
wire signed[31:0]    reg_psum_28_9;
wire signed[31:0]    reg_weight_28_10;
wire signed[31:0]    reg_psum_28_10;
wire signed[31:0]    reg_weight_28_11;
wire signed[31:0]    reg_psum_28_11;
wire signed[31:0]    reg_weight_28_12;
wire signed[31:0]    reg_psum_28_12;
wire signed[31:0]    reg_weight_28_13;
wire signed[31:0]    reg_psum_28_13;
wire signed[31:0]    reg_weight_28_14;
wire signed[31:0]    reg_psum_28_14;
wire signed[31:0]    reg_weight_28_15;
wire signed[31:0]    reg_psum_28_15;
wire signed[31:0]    reg_weight_28_16;
wire signed[31:0]    reg_psum_28_16;
wire signed[31:0]    reg_weight_28_17;
wire signed[31:0]    reg_psum_28_17;
wire signed[31:0]    reg_weight_28_18;
wire signed[31:0]    reg_psum_28_18;
wire signed[31:0]    reg_weight_28_19;
wire signed[31:0]    reg_psum_28_19;
wire signed[31:0]    reg_weight_28_20;
wire signed[31:0]    reg_psum_28_20;
wire signed[31:0]    reg_weight_28_21;
wire signed[31:0]    reg_psum_28_21;
wire signed[31:0]    reg_weight_28_22;
wire signed[31:0]    reg_psum_28_22;
wire signed[31:0]    reg_weight_28_23;
wire signed[31:0]    reg_psum_28_23;
wire signed[31:0]    reg_weight_28_24;
wire signed[31:0]    reg_psum_28_24;
wire signed[31:0]    reg_weight_28_25;
wire signed[31:0]    reg_psum_28_25;
wire signed[31:0]    reg_weight_28_26;
wire signed[31:0]    reg_psum_28_26;
wire signed[31:0]    reg_weight_28_27;
wire signed[31:0]    reg_psum_28_27;
wire signed[31:0]    reg_weight_28_28;
wire signed[31:0]    reg_psum_28_28;
wire signed[31:0]    reg_weight_28_29;
wire signed[31:0]    reg_psum_28_29;
wire signed[31:0]    reg_weight_28_30;
wire signed[31:0]    reg_psum_28_30;
wire signed[31:0]    reg_weight_28_31;
wire signed[31:0]    reg_psum_28_31;
wire signed[31:0]    reg_weight_28_32;
wire signed[31:0]    reg_psum_28_32;
wire signed[31:0]    reg_weight_28_33;
wire signed[31:0]    reg_psum_28_33;
wire signed[31:0]    reg_weight_28_34;
wire signed[31:0]    reg_psum_28_34;
wire signed[31:0]    reg_weight_28_35;
wire signed[31:0]    reg_psum_28_35;
wire signed[31:0]    reg_weight_28_36;
wire signed[31:0]    reg_psum_28_36;
wire signed[31:0]    reg_weight_28_37;
wire signed[31:0]    reg_psum_28_37;
wire signed[31:0]    reg_weight_28_38;
wire signed[31:0]    reg_psum_28_38;
wire signed[31:0]    reg_weight_28_39;
wire signed[31:0]    reg_psum_28_39;
wire signed[31:0]    reg_weight_28_40;
wire signed[31:0]    reg_psum_28_40;
wire signed[31:0]    reg_weight_28_41;
wire signed[31:0]    reg_psum_28_41;
wire signed[31:0]    reg_weight_28_42;
wire signed[31:0]    reg_psum_28_42;
wire signed[31:0]    reg_weight_28_43;
wire signed[31:0]    reg_psum_28_43;
wire signed[31:0]    reg_weight_28_44;
wire signed[31:0]    reg_psum_28_44;
wire signed[31:0]    reg_weight_28_45;
wire signed[31:0]    reg_psum_28_45;
wire signed[31:0]    reg_weight_28_46;
wire signed[31:0]    reg_psum_28_46;
wire signed[31:0]    reg_weight_28_47;
wire signed[31:0]    reg_psum_28_47;
wire signed[31:0]    reg_weight_28_48;
wire signed[31:0]    reg_psum_28_48;
wire signed[31:0]    reg_weight_28_49;
wire signed[31:0]    reg_psum_28_49;
wire signed[31:0]    reg_weight_28_50;
wire signed[31:0]    reg_psum_28_50;
wire signed[31:0]    reg_weight_28_51;
wire signed[31:0]    reg_psum_28_51;
wire signed[31:0]    reg_weight_28_52;
wire signed[31:0]    reg_psum_28_52;
wire signed[31:0]    reg_weight_28_53;
wire signed[31:0]    reg_psum_28_53;
wire signed[31:0]    reg_weight_28_54;
wire signed[31:0]    reg_psum_28_54;
wire signed[31:0]    reg_weight_28_55;
wire signed[31:0]    reg_psum_28_55;
wire signed[31:0]    reg_weight_28_56;
wire signed[31:0]    reg_psum_28_56;
wire signed[31:0]    reg_weight_28_57;
wire signed[31:0]    reg_psum_28_57;
wire signed[31:0]    reg_weight_28_58;
wire signed[31:0]    reg_psum_28_58;
wire signed[31:0]    reg_weight_28_59;
wire signed[31:0]    reg_psum_28_59;
wire signed[31:0]    reg_weight_28_60;
wire signed[31:0]    reg_psum_28_60;
wire signed[31:0]    reg_weight_28_61;
wire signed[31:0]    reg_psum_28_61;
wire signed[31:0]    reg_weight_28_62;
wire signed[31:0]    reg_psum_28_62;
wire signed[31:0]    reg_weight_28_63;
wire signed[31:0]    reg_psum_28_63;
wire signed[31:0]    reg_weight_29_0;
wire signed[31:0]    reg_psum_29_0;
wire signed[31:0]    reg_weight_29_1;
wire signed[31:0]    reg_psum_29_1;
wire signed[31:0]    reg_weight_29_2;
wire signed[31:0]    reg_psum_29_2;
wire signed[31:0]    reg_weight_29_3;
wire signed[31:0]    reg_psum_29_3;
wire signed[31:0]    reg_weight_29_4;
wire signed[31:0]    reg_psum_29_4;
wire signed[31:0]    reg_weight_29_5;
wire signed[31:0]    reg_psum_29_5;
wire signed[31:0]    reg_weight_29_6;
wire signed[31:0]    reg_psum_29_6;
wire signed[31:0]    reg_weight_29_7;
wire signed[31:0]    reg_psum_29_7;
wire signed[31:0]    reg_weight_29_8;
wire signed[31:0]    reg_psum_29_8;
wire signed[31:0]    reg_weight_29_9;
wire signed[31:0]    reg_psum_29_9;
wire signed[31:0]    reg_weight_29_10;
wire signed[31:0]    reg_psum_29_10;
wire signed[31:0]    reg_weight_29_11;
wire signed[31:0]    reg_psum_29_11;
wire signed[31:0]    reg_weight_29_12;
wire signed[31:0]    reg_psum_29_12;
wire signed[31:0]    reg_weight_29_13;
wire signed[31:0]    reg_psum_29_13;
wire signed[31:0]    reg_weight_29_14;
wire signed[31:0]    reg_psum_29_14;
wire signed[31:0]    reg_weight_29_15;
wire signed[31:0]    reg_psum_29_15;
wire signed[31:0]    reg_weight_29_16;
wire signed[31:0]    reg_psum_29_16;
wire signed[31:0]    reg_weight_29_17;
wire signed[31:0]    reg_psum_29_17;
wire signed[31:0]    reg_weight_29_18;
wire signed[31:0]    reg_psum_29_18;
wire signed[31:0]    reg_weight_29_19;
wire signed[31:0]    reg_psum_29_19;
wire signed[31:0]    reg_weight_29_20;
wire signed[31:0]    reg_psum_29_20;
wire signed[31:0]    reg_weight_29_21;
wire signed[31:0]    reg_psum_29_21;
wire signed[31:0]    reg_weight_29_22;
wire signed[31:0]    reg_psum_29_22;
wire signed[31:0]    reg_weight_29_23;
wire signed[31:0]    reg_psum_29_23;
wire signed[31:0]    reg_weight_29_24;
wire signed[31:0]    reg_psum_29_24;
wire signed[31:0]    reg_weight_29_25;
wire signed[31:0]    reg_psum_29_25;
wire signed[31:0]    reg_weight_29_26;
wire signed[31:0]    reg_psum_29_26;
wire signed[31:0]    reg_weight_29_27;
wire signed[31:0]    reg_psum_29_27;
wire signed[31:0]    reg_weight_29_28;
wire signed[31:0]    reg_psum_29_28;
wire signed[31:0]    reg_weight_29_29;
wire signed[31:0]    reg_psum_29_29;
wire signed[31:0]    reg_weight_29_30;
wire signed[31:0]    reg_psum_29_30;
wire signed[31:0]    reg_weight_29_31;
wire signed[31:0]    reg_psum_29_31;
wire signed[31:0]    reg_weight_29_32;
wire signed[31:0]    reg_psum_29_32;
wire signed[31:0]    reg_weight_29_33;
wire signed[31:0]    reg_psum_29_33;
wire signed[31:0]    reg_weight_29_34;
wire signed[31:0]    reg_psum_29_34;
wire signed[31:0]    reg_weight_29_35;
wire signed[31:0]    reg_psum_29_35;
wire signed[31:0]    reg_weight_29_36;
wire signed[31:0]    reg_psum_29_36;
wire signed[31:0]    reg_weight_29_37;
wire signed[31:0]    reg_psum_29_37;
wire signed[31:0]    reg_weight_29_38;
wire signed[31:0]    reg_psum_29_38;
wire signed[31:0]    reg_weight_29_39;
wire signed[31:0]    reg_psum_29_39;
wire signed[31:0]    reg_weight_29_40;
wire signed[31:0]    reg_psum_29_40;
wire signed[31:0]    reg_weight_29_41;
wire signed[31:0]    reg_psum_29_41;
wire signed[31:0]    reg_weight_29_42;
wire signed[31:0]    reg_psum_29_42;
wire signed[31:0]    reg_weight_29_43;
wire signed[31:0]    reg_psum_29_43;
wire signed[31:0]    reg_weight_29_44;
wire signed[31:0]    reg_psum_29_44;
wire signed[31:0]    reg_weight_29_45;
wire signed[31:0]    reg_psum_29_45;
wire signed[31:0]    reg_weight_29_46;
wire signed[31:0]    reg_psum_29_46;
wire signed[31:0]    reg_weight_29_47;
wire signed[31:0]    reg_psum_29_47;
wire signed[31:0]    reg_weight_29_48;
wire signed[31:0]    reg_psum_29_48;
wire signed[31:0]    reg_weight_29_49;
wire signed[31:0]    reg_psum_29_49;
wire signed[31:0]    reg_weight_29_50;
wire signed[31:0]    reg_psum_29_50;
wire signed[31:0]    reg_weight_29_51;
wire signed[31:0]    reg_psum_29_51;
wire signed[31:0]    reg_weight_29_52;
wire signed[31:0]    reg_psum_29_52;
wire signed[31:0]    reg_weight_29_53;
wire signed[31:0]    reg_psum_29_53;
wire signed[31:0]    reg_weight_29_54;
wire signed[31:0]    reg_psum_29_54;
wire signed[31:0]    reg_weight_29_55;
wire signed[31:0]    reg_psum_29_55;
wire signed[31:0]    reg_weight_29_56;
wire signed[31:0]    reg_psum_29_56;
wire signed[31:0]    reg_weight_29_57;
wire signed[31:0]    reg_psum_29_57;
wire signed[31:0]    reg_weight_29_58;
wire signed[31:0]    reg_psum_29_58;
wire signed[31:0]    reg_weight_29_59;
wire signed[31:0]    reg_psum_29_59;
wire signed[31:0]    reg_weight_29_60;
wire signed[31:0]    reg_psum_29_60;
wire signed[31:0]    reg_weight_29_61;
wire signed[31:0]    reg_psum_29_61;
wire signed[31:0]    reg_weight_29_62;
wire signed[31:0]    reg_psum_29_62;
wire signed[31:0]    reg_weight_29_63;
wire signed[31:0]    reg_psum_29_63;
wire signed[31:0]    reg_weight_30_0;
wire signed[31:0]    reg_psum_30_0;
wire signed[31:0]    reg_weight_30_1;
wire signed[31:0]    reg_psum_30_1;
wire signed[31:0]    reg_weight_30_2;
wire signed[31:0]    reg_psum_30_2;
wire signed[31:0]    reg_weight_30_3;
wire signed[31:0]    reg_psum_30_3;
wire signed[31:0]    reg_weight_30_4;
wire signed[31:0]    reg_psum_30_4;
wire signed[31:0]    reg_weight_30_5;
wire signed[31:0]    reg_psum_30_5;
wire signed[31:0]    reg_weight_30_6;
wire signed[31:0]    reg_psum_30_6;
wire signed[31:0]    reg_weight_30_7;
wire signed[31:0]    reg_psum_30_7;
wire signed[31:0]    reg_weight_30_8;
wire signed[31:0]    reg_psum_30_8;
wire signed[31:0]    reg_weight_30_9;
wire signed[31:0]    reg_psum_30_9;
wire signed[31:0]    reg_weight_30_10;
wire signed[31:0]    reg_psum_30_10;
wire signed[31:0]    reg_weight_30_11;
wire signed[31:0]    reg_psum_30_11;
wire signed[31:0]    reg_weight_30_12;
wire signed[31:0]    reg_psum_30_12;
wire signed[31:0]    reg_weight_30_13;
wire signed[31:0]    reg_psum_30_13;
wire signed[31:0]    reg_weight_30_14;
wire signed[31:0]    reg_psum_30_14;
wire signed[31:0]    reg_weight_30_15;
wire signed[31:0]    reg_psum_30_15;
wire signed[31:0]    reg_weight_30_16;
wire signed[31:0]    reg_psum_30_16;
wire signed[31:0]    reg_weight_30_17;
wire signed[31:0]    reg_psum_30_17;
wire signed[31:0]    reg_weight_30_18;
wire signed[31:0]    reg_psum_30_18;
wire signed[31:0]    reg_weight_30_19;
wire signed[31:0]    reg_psum_30_19;
wire signed[31:0]    reg_weight_30_20;
wire signed[31:0]    reg_psum_30_20;
wire signed[31:0]    reg_weight_30_21;
wire signed[31:0]    reg_psum_30_21;
wire signed[31:0]    reg_weight_30_22;
wire signed[31:0]    reg_psum_30_22;
wire signed[31:0]    reg_weight_30_23;
wire signed[31:0]    reg_psum_30_23;
wire signed[31:0]    reg_weight_30_24;
wire signed[31:0]    reg_psum_30_24;
wire signed[31:0]    reg_weight_30_25;
wire signed[31:0]    reg_psum_30_25;
wire signed[31:0]    reg_weight_30_26;
wire signed[31:0]    reg_psum_30_26;
wire signed[31:0]    reg_weight_30_27;
wire signed[31:0]    reg_psum_30_27;
wire signed[31:0]    reg_weight_30_28;
wire signed[31:0]    reg_psum_30_28;
wire signed[31:0]    reg_weight_30_29;
wire signed[31:0]    reg_psum_30_29;
wire signed[31:0]    reg_weight_30_30;
wire signed[31:0]    reg_psum_30_30;
wire signed[31:0]    reg_weight_30_31;
wire signed[31:0]    reg_psum_30_31;
wire signed[31:0]    reg_weight_30_32;
wire signed[31:0]    reg_psum_30_32;
wire signed[31:0]    reg_weight_30_33;
wire signed[31:0]    reg_psum_30_33;
wire signed[31:0]    reg_weight_30_34;
wire signed[31:0]    reg_psum_30_34;
wire signed[31:0]    reg_weight_30_35;
wire signed[31:0]    reg_psum_30_35;
wire signed[31:0]    reg_weight_30_36;
wire signed[31:0]    reg_psum_30_36;
wire signed[31:0]    reg_weight_30_37;
wire signed[31:0]    reg_psum_30_37;
wire signed[31:0]    reg_weight_30_38;
wire signed[31:0]    reg_psum_30_38;
wire signed[31:0]    reg_weight_30_39;
wire signed[31:0]    reg_psum_30_39;
wire signed[31:0]    reg_weight_30_40;
wire signed[31:0]    reg_psum_30_40;
wire signed[31:0]    reg_weight_30_41;
wire signed[31:0]    reg_psum_30_41;
wire signed[31:0]    reg_weight_30_42;
wire signed[31:0]    reg_psum_30_42;
wire signed[31:0]    reg_weight_30_43;
wire signed[31:0]    reg_psum_30_43;
wire signed[31:0]    reg_weight_30_44;
wire signed[31:0]    reg_psum_30_44;
wire signed[31:0]    reg_weight_30_45;
wire signed[31:0]    reg_psum_30_45;
wire signed[31:0]    reg_weight_30_46;
wire signed[31:0]    reg_psum_30_46;
wire signed[31:0]    reg_weight_30_47;
wire signed[31:0]    reg_psum_30_47;
wire signed[31:0]    reg_weight_30_48;
wire signed[31:0]    reg_psum_30_48;
wire signed[31:0]    reg_weight_30_49;
wire signed[31:0]    reg_psum_30_49;
wire signed[31:0]    reg_weight_30_50;
wire signed[31:0]    reg_psum_30_50;
wire signed[31:0]    reg_weight_30_51;
wire signed[31:0]    reg_psum_30_51;
wire signed[31:0]    reg_weight_30_52;
wire signed[31:0]    reg_psum_30_52;
wire signed[31:0]    reg_weight_30_53;
wire signed[31:0]    reg_psum_30_53;
wire signed[31:0]    reg_weight_30_54;
wire signed[31:0]    reg_psum_30_54;
wire signed[31:0]    reg_weight_30_55;
wire signed[31:0]    reg_psum_30_55;
wire signed[31:0]    reg_weight_30_56;
wire signed[31:0]    reg_psum_30_56;
wire signed[31:0]    reg_weight_30_57;
wire signed[31:0]    reg_psum_30_57;
wire signed[31:0]    reg_weight_30_58;
wire signed[31:0]    reg_psum_30_58;
wire signed[31:0]    reg_weight_30_59;
wire signed[31:0]    reg_psum_30_59;
wire signed[31:0]    reg_weight_30_60;
wire signed[31:0]    reg_psum_30_60;
wire signed[31:0]    reg_weight_30_61;
wire signed[31:0]    reg_psum_30_61;
wire signed[31:0]    reg_weight_30_62;
wire signed[31:0]    reg_psum_30_62;
wire signed[31:0]    reg_weight_30_63;
wire signed[31:0]    reg_psum_30_63;
wire signed[31:0]    reg_weight_31_0;
wire signed[31:0]    reg_psum_31_0;
wire signed[31:0]    reg_weight_31_1;
wire signed[31:0]    reg_psum_31_1;
wire signed[31:0]    reg_weight_31_2;
wire signed[31:0]    reg_psum_31_2;
wire signed[31:0]    reg_weight_31_3;
wire signed[31:0]    reg_psum_31_3;
wire signed[31:0]    reg_weight_31_4;
wire signed[31:0]    reg_psum_31_4;
wire signed[31:0]    reg_weight_31_5;
wire signed[31:0]    reg_psum_31_5;
wire signed[31:0]    reg_weight_31_6;
wire signed[31:0]    reg_psum_31_6;
wire signed[31:0]    reg_weight_31_7;
wire signed[31:0]    reg_psum_31_7;
wire signed[31:0]    reg_weight_31_8;
wire signed[31:0]    reg_psum_31_8;
wire signed[31:0]    reg_weight_31_9;
wire signed[31:0]    reg_psum_31_9;
wire signed[31:0]    reg_weight_31_10;
wire signed[31:0]    reg_psum_31_10;
wire signed[31:0]    reg_weight_31_11;
wire signed[31:0]    reg_psum_31_11;
wire signed[31:0]    reg_weight_31_12;
wire signed[31:0]    reg_psum_31_12;
wire signed[31:0]    reg_weight_31_13;
wire signed[31:0]    reg_psum_31_13;
wire signed[31:0]    reg_weight_31_14;
wire signed[31:0]    reg_psum_31_14;
wire signed[31:0]    reg_weight_31_15;
wire signed[31:0]    reg_psum_31_15;
wire signed[31:0]    reg_weight_31_16;
wire signed[31:0]    reg_psum_31_16;
wire signed[31:0]    reg_weight_31_17;
wire signed[31:0]    reg_psum_31_17;
wire signed[31:0]    reg_weight_31_18;
wire signed[31:0]    reg_psum_31_18;
wire signed[31:0]    reg_weight_31_19;
wire signed[31:0]    reg_psum_31_19;
wire signed[31:0]    reg_weight_31_20;
wire signed[31:0]    reg_psum_31_20;
wire signed[31:0]    reg_weight_31_21;
wire signed[31:0]    reg_psum_31_21;
wire signed[31:0]    reg_weight_31_22;
wire signed[31:0]    reg_psum_31_22;
wire signed[31:0]    reg_weight_31_23;
wire signed[31:0]    reg_psum_31_23;
wire signed[31:0]    reg_weight_31_24;
wire signed[31:0]    reg_psum_31_24;
wire signed[31:0]    reg_weight_31_25;
wire signed[31:0]    reg_psum_31_25;
wire signed[31:0]    reg_weight_31_26;
wire signed[31:0]    reg_psum_31_26;
wire signed[31:0]    reg_weight_31_27;
wire signed[31:0]    reg_psum_31_27;
wire signed[31:0]    reg_weight_31_28;
wire signed[31:0]    reg_psum_31_28;
wire signed[31:0]    reg_weight_31_29;
wire signed[31:0]    reg_psum_31_29;
wire signed[31:0]    reg_weight_31_30;
wire signed[31:0]    reg_psum_31_30;
wire signed[31:0]    reg_weight_31_31;
wire signed[31:0]    reg_psum_31_31;
wire signed[31:0]    reg_weight_31_32;
wire signed[31:0]    reg_psum_31_32;
wire signed[31:0]    reg_weight_31_33;
wire signed[31:0]    reg_psum_31_33;
wire signed[31:0]    reg_weight_31_34;
wire signed[31:0]    reg_psum_31_34;
wire signed[31:0]    reg_weight_31_35;
wire signed[31:0]    reg_psum_31_35;
wire signed[31:0]    reg_weight_31_36;
wire signed[31:0]    reg_psum_31_36;
wire signed[31:0]    reg_weight_31_37;
wire signed[31:0]    reg_psum_31_37;
wire signed[31:0]    reg_weight_31_38;
wire signed[31:0]    reg_psum_31_38;
wire signed[31:0]    reg_weight_31_39;
wire signed[31:0]    reg_psum_31_39;
wire signed[31:0]    reg_weight_31_40;
wire signed[31:0]    reg_psum_31_40;
wire signed[31:0]    reg_weight_31_41;
wire signed[31:0]    reg_psum_31_41;
wire signed[31:0]    reg_weight_31_42;
wire signed[31:0]    reg_psum_31_42;
wire signed[31:0]    reg_weight_31_43;
wire signed[31:0]    reg_psum_31_43;
wire signed[31:0]    reg_weight_31_44;
wire signed[31:0]    reg_psum_31_44;
wire signed[31:0]    reg_weight_31_45;
wire signed[31:0]    reg_psum_31_45;
wire signed[31:0]    reg_weight_31_46;
wire signed[31:0]    reg_psum_31_46;
wire signed[31:0]    reg_weight_31_47;
wire signed[31:0]    reg_psum_31_47;
wire signed[31:0]    reg_weight_31_48;
wire signed[31:0]    reg_psum_31_48;
wire signed[31:0]    reg_weight_31_49;
wire signed[31:0]    reg_psum_31_49;
wire signed[31:0]    reg_weight_31_50;
wire signed[31:0]    reg_psum_31_50;
wire signed[31:0]    reg_weight_31_51;
wire signed[31:0]    reg_psum_31_51;
wire signed[31:0]    reg_weight_31_52;
wire signed[31:0]    reg_psum_31_52;
wire signed[31:0]    reg_weight_31_53;
wire signed[31:0]    reg_psum_31_53;
wire signed[31:0]    reg_weight_31_54;
wire signed[31:0]    reg_psum_31_54;
wire signed[31:0]    reg_weight_31_55;
wire signed[31:0]    reg_psum_31_55;
wire signed[31:0]    reg_weight_31_56;
wire signed[31:0]    reg_psum_31_56;
wire signed[31:0]    reg_weight_31_57;
wire signed[31:0]    reg_psum_31_57;
wire signed[31:0]    reg_weight_31_58;
wire signed[31:0]    reg_psum_31_58;
wire signed[31:0]    reg_weight_31_59;
wire signed[31:0]    reg_psum_31_59;
wire signed[31:0]    reg_weight_31_60;
wire signed[31:0]    reg_psum_31_60;
wire signed[31:0]    reg_weight_31_61;
wire signed[31:0]    reg_psum_31_61;
wire signed[31:0]    reg_weight_31_62;
wire signed[31:0]    reg_psum_31_62;
wire signed[31:0]    reg_weight_31_63;
wire signed[31:0]    reg_psum_31_63;
wire signed[31:0]    reg_weight_32_0;
wire signed[31:0]    reg_psum_32_0;
wire signed[31:0]    reg_weight_32_1;
wire signed[31:0]    reg_psum_32_1;
wire signed[31:0]    reg_weight_32_2;
wire signed[31:0]    reg_psum_32_2;
wire signed[31:0]    reg_weight_32_3;
wire signed[31:0]    reg_psum_32_3;
wire signed[31:0]    reg_weight_32_4;
wire signed[31:0]    reg_psum_32_4;
wire signed[31:0]    reg_weight_32_5;
wire signed[31:0]    reg_psum_32_5;
wire signed[31:0]    reg_weight_32_6;
wire signed[31:0]    reg_psum_32_6;
wire signed[31:0]    reg_weight_32_7;
wire signed[31:0]    reg_psum_32_7;
wire signed[31:0]    reg_weight_32_8;
wire signed[31:0]    reg_psum_32_8;
wire signed[31:0]    reg_weight_32_9;
wire signed[31:0]    reg_psum_32_9;
wire signed[31:0]    reg_weight_32_10;
wire signed[31:0]    reg_psum_32_10;
wire signed[31:0]    reg_weight_32_11;
wire signed[31:0]    reg_psum_32_11;
wire signed[31:0]    reg_weight_32_12;
wire signed[31:0]    reg_psum_32_12;
wire signed[31:0]    reg_weight_32_13;
wire signed[31:0]    reg_psum_32_13;
wire signed[31:0]    reg_weight_32_14;
wire signed[31:0]    reg_psum_32_14;
wire signed[31:0]    reg_weight_32_15;
wire signed[31:0]    reg_psum_32_15;
wire signed[31:0]    reg_weight_32_16;
wire signed[31:0]    reg_psum_32_16;
wire signed[31:0]    reg_weight_32_17;
wire signed[31:0]    reg_psum_32_17;
wire signed[31:0]    reg_weight_32_18;
wire signed[31:0]    reg_psum_32_18;
wire signed[31:0]    reg_weight_32_19;
wire signed[31:0]    reg_psum_32_19;
wire signed[31:0]    reg_weight_32_20;
wire signed[31:0]    reg_psum_32_20;
wire signed[31:0]    reg_weight_32_21;
wire signed[31:0]    reg_psum_32_21;
wire signed[31:0]    reg_weight_32_22;
wire signed[31:0]    reg_psum_32_22;
wire signed[31:0]    reg_weight_32_23;
wire signed[31:0]    reg_psum_32_23;
wire signed[31:0]    reg_weight_32_24;
wire signed[31:0]    reg_psum_32_24;
wire signed[31:0]    reg_weight_32_25;
wire signed[31:0]    reg_psum_32_25;
wire signed[31:0]    reg_weight_32_26;
wire signed[31:0]    reg_psum_32_26;
wire signed[31:0]    reg_weight_32_27;
wire signed[31:0]    reg_psum_32_27;
wire signed[31:0]    reg_weight_32_28;
wire signed[31:0]    reg_psum_32_28;
wire signed[31:0]    reg_weight_32_29;
wire signed[31:0]    reg_psum_32_29;
wire signed[31:0]    reg_weight_32_30;
wire signed[31:0]    reg_psum_32_30;
wire signed[31:0]    reg_weight_32_31;
wire signed[31:0]    reg_psum_32_31;
wire signed[31:0]    reg_weight_32_32;
wire signed[31:0]    reg_psum_32_32;
wire signed[31:0]    reg_weight_32_33;
wire signed[31:0]    reg_psum_32_33;
wire signed[31:0]    reg_weight_32_34;
wire signed[31:0]    reg_psum_32_34;
wire signed[31:0]    reg_weight_32_35;
wire signed[31:0]    reg_psum_32_35;
wire signed[31:0]    reg_weight_32_36;
wire signed[31:0]    reg_psum_32_36;
wire signed[31:0]    reg_weight_32_37;
wire signed[31:0]    reg_psum_32_37;
wire signed[31:0]    reg_weight_32_38;
wire signed[31:0]    reg_psum_32_38;
wire signed[31:0]    reg_weight_32_39;
wire signed[31:0]    reg_psum_32_39;
wire signed[31:0]    reg_weight_32_40;
wire signed[31:0]    reg_psum_32_40;
wire signed[31:0]    reg_weight_32_41;
wire signed[31:0]    reg_psum_32_41;
wire signed[31:0]    reg_weight_32_42;
wire signed[31:0]    reg_psum_32_42;
wire signed[31:0]    reg_weight_32_43;
wire signed[31:0]    reg_psum_32_43;
wire signed[31:0]    reg_weight_32_44;
wire signed[31:0]    reg_psum_32_44;
wire signed[31:0]    reg_weight_32_45;
wire signed[31:0]    reg_psum_32_45;
wire signed[31:0]    reg_weight_32_46;
wire signed[31:0]    reg_psum_32_46;
wire signed[31:0]    reg_weight_32_47;
wire signed[31:0]    reg_psum_32_47;
wire signed[31:0]    reg_weight_32_48;
wire signed[31:0]    reg_psum_32_48;
wire signed[31:0]    reg_weight_32_49;
wire signed[31:0]    reg_psum_32_49;
wire signed[31:0]    reg_weight_32_50;
wire signed[31:0]    reg_psum_32_50;
wire signed[31:0]    reg_weight_32_51;
wire signed[31:0]    reg_psum_32_51;
wire signed[31:0]    reg_weight_32_52;
wire signed[31:0]    reg_psum_32_52;
wire signed[31:0]    reg_weight_32_53;
wire signed[31:0]    reg_psum_32_53;
wire signed[31:0]    reg_weight_32_54;
wire signed[31:0]    reg_psum_32_54;
wire signed[31:0]    reg_weight_32_55;
wire signed[31:0]    reg_psum_32_55;
wire signed[31:0]    reg_weight_32_56;
wire signed[31:0]    reg_psum_32_56;
wire signed[31:0]    reg_weight_32_57;
wire signed[31:0]    reg_psum_32_57;
wire signed[31:0]    reg_weight_32_58;
wire signed[31:0]    reg_psum_32_58;
wire signed[31:0]    reg_weight_32_59;
wire signed[31:0]    reg_psum_32_59;
wire signed[31:0]    reg_weight_32_60;
wire signed[31:0]    reg_psum_32_60;
wire signed[31:0]    reg_weight_32_61;
wire signed[31:0]    reg_psum_32_61;
wire signed[31:0]    reg_weight_32_62;
wire signed[31:0]    reg_psum_32_62;
wire signed[31:0]    reg_weight_32_63;
wire signed[31:0]    reg_psum_32_63;
wire signed[31:0]    reg_weight_33_0;
wire signed[31:0]    reg_psum_33_0;
wire signed[31:0]    reg_weight_33_1;
wire signed[31:0]    reg_psum_33_1;
wire signed[31:0]    reg_weight_33_2;
wire signed[31:0]    reg_psum_33_2;
wire signed[31:0]    reg_weight_33_3;
wire signed[31:0]    reg_psum_33_3;
wire signed[31:0]    reg_weight_33_4;
wire signed[31:0]    reg_psum_33_4;
wire signed[31:0]    reg_weight_33_5;
wire signed[31:0]    reg_psum_33_5;
wire signed[31:0]    reg_weight_33_6;
wire signed[31:0]    reg_psum_33_6;
wire signed[31:0]    reg_weight_33_7;
wire signed[31:0]    reg_psum_33_7;
wire signed[31:0]    reg_weight_33_8;
wire signed[31:0]    reg_psum_33_8;
wire signed[31:0]    reg_weight_33_9;
wire signed[31:0]    reg_psum_33_9;
wire signed[31:0]    reg_weight_33_10;
wire signed[31:0]    reg_psum_33_10;
wire signed[31:0]    reg_weight_33_11;
wire signed[31:0]    reg_psum_33_11;
wire signed[31:0]    reg_weight_33_12;
wire signed[31:0]    reg_psum_33_12;
wire signed[31:0]    reg_weight_33_13;
wire signed[31:0]    reg_psum_33_13;
wire signed[31:0]    reg_weight_33_14;
wire signed[31:0]    reg_psum_33_14;
wire signed[31:0]    reg_weight_33_15;
wire signed[31:0]    reg_psum_33_15;
wire signed[31:0]    reg_weight_33_16;
wire signed[31:0]    reg_psum_33_16;
wire signed[31:0]    reg_weight_33_17;
wire signed[31:0]    reg_psum_33_17;
wire signed[31:0]    reg_weight_33_18;
wire signed[31:0]    reg_psum_33_18;
wire signed[31:0]    reg_weight_33_19;
wire signed[31:0]    reg_psum_33_19;
wire signed[31:0]    reg_weight_33_20;
wire signed[31:0]    reg_psum_33_20;
wire signed[31:0]    reg_weight_33_21;
wire signed[31:0]    reg_psum_33_21;
wire signed[31:0]    reg_weight_33_22;
wire signed[31:0]    reg_psum_33_22;
wire signed[31:0]    reg_weight_33_23;
wire signed[31:0]    reg_psum_33_23;
wire signed[31:0]    reg_weight_33_24;
wire signed[31:0]    reg_psum_33_24;
wire signed[31:0]    reg_weight_33_25;
wire signed[31:0]    reg_psum_33_25;
wire signed[31:0]    reg_weight_33_26;
wire signed[31:0]    reg_psum_33_26;
wire signed[31:0]    reg_weight_33_27;
wire signed[31:0]    reg_psum_33_27;
wire signed[31:0]    reg_weight_33_28;
wire signed[31:0]    reg_psum_33_28;
wire signed[31:0]    reg_weight_33_29;
wire signed[31:0]    reg_psum_33_29;
wire signed[31:0]    reg_weight_33_30;
wire signed[31:0]    reg_psum_33_30;
wire signed[31:0]    reg_weight_33_31;
wire signed[31:0]    reg_psum_33_31;
wire signed[31:0]    reg_weight_33_32;
wire signed[31:0]    reg_psum_33_32;
wire signed[31:0]    reg_weight_33_33;
wire signed[31:0]    reg_psum_33_33;
wire signed[31:0]    reg_weight_33_34;
wire signed[31:0]    reg_psum_33_34;
wire signed[31:0]    reg_weight_33_35;
wire signed[31:0]    reg_psum_33_35;
wire signed[31:0]    reg_weight_33_36;
wire signed[31:0]    reg_psum_33_36;
wire signed[31:0]    reg_weight_33_37;
wire signed[31:0]    reg_psum_33_37;
wire signed[31:0]    reg_weight_33_38;
wire signed[31:0]    reg_psum_33_38;
wire signed[31:0]    reg_weight_33_39;
wire signed[31:0]    reg_psum_33_39;
wire signed[31:0]    reg_weight_33_40;
wire signed[31:0]    reg_psum_33_40;
wire signed[31:0]    reg_weight_33_41;
wire signed[31:0]    reg_psum_33_41;
wire signed[31:0]    reg_weight_33_42;
wire signed[31:0]    reg_psum_33_42;
wire signed[31:0]    reg_weight_33_43;
wire signed[31:0]    reg_psum_33_43;
wire signed[31:0]    reg_weight_33_44;
wire signed[31:0]    reg_psum_33_44;
wire signed[31:0]    reg_weight_33_45;
wire signed[31:0]    reg_psum_33_45;
wire signed[31:0]    reg_weight_33_46;
wire signed[31:0]    reg_psum_33_46;
wire signed[31:0]    reg_weight_33_47;
wire signed[31:0]    reg_psum_33_47;
wire signed[31:0]    reg_weight_33_48;
wire signed[31:0]    reg_psum_33_48;
wire signed[31:0]    reg_weight_33_49;
wire signed[31:0]    reg_psum_33_49;
wire signed[31:0]    reg_weight_33_50;
wire signed[31:0]    reg_psum_33_50;
wire signed[31:0]    reg_weight_33_51;
wire signed[31:0]    reg_psum_33_51;
wire signed[31:0]    reg_weight_33_52;
wire signed[31:0]    reg_psum_33_52;
wire signed[31:0]    reg_weight_33_53;
wire signed[31:0]    reg_psum_33_53;
wire signed[31:0]    reg_weight_33_54;
wire signed[31:0]    reg_psum_33_54;
wire signed[31:0]    reg_weight_33_55;
wire signed[31:0]    reg_psum_33_55;
wire signed[31:0]    reg_weight_33_56;
wire signed[31:0]    reg_psum_33_56;
wire signed[31:0]    reg_weight_33_57;
wire signed[31:0]    reg_psum_33_57;
wire signed[31:0]    reg_weight_33_58;
wire signed[31:0]    reg_psum_33_58;
wire signed[31:0]    reg_weight_33_59;
wire signed[31:0]    reg_psum_33_59;
wire signed[31:0]    reg_weight_33_60;
wire signed[31:0]    reg_psum_33_60;
wire signed[31:0]    reg_weight_33_61;
wire signed[31:0]    reg_psum_33_61;
wire signed[31:0]    reg_weight_33_62;
wire signed[31:0]    reg_psum_33_62;
wire signed[31:0]    reg_weight_33_63;
wire signed[31:0]    reg_psum_33_63;
wire signed[31:0]    reg_weight_34_0;
wire signed[31:0]    reg_psum_34_0;
wire signed[31:0]    reg_weight_34_1;
wire signed[31:0]    reg_psum_34_1;
wire signed[31:0]    reg_weight_34_2;
wire signed[31:0]    reg_psum_34_2;
wire signed[31:0]    reg_weight_34_3;
wire signed[31:0]    reg_psum_34_3;
wire signed[31:0]    reg_weight_34_4;
wire signed[31:0]    reg_psum_34_4;
wire signed[31:0]    reg_weight_34_5;
wire signed[31:0]    reg_psum_34_5;
wire signed[31:0]    reg_weight_34_6;
wire signed[31:0]    reg_psum_34_6;
wire signed[31:0]    reg_weight_34_7;
wire signed[31:0]    reg_psum_34_7;
wire signed[31:0]    reg_weight_34_8;
wire signed[31:0]    reg_psum_34_8;
wire signed[31:0]    reg_weight_34_9;
wire signed[31:0]    reg_psum_34_9;
wire signed[31:0]    reg_weight_34_10;
wire signed[31:0]    reg_psum_34_10;
wire signed[31:0]    reg_weight_34_11;
wire signed[31:0]    reg_psum_34_11;
wire signed[31:0]    reg_weight_34_12;
wire signed[31:0]    reg_psum_34_12;
wire signed[31:0]    reg_weight_34_13;
wire signed[31:0]    reg_psum_34_13;
wire signed[31:0]    reg_weight_34_14;
wire signed[31:0]    reg_psum_34_14;
wire signed[31:0]    reg_weight_34_15;
wire signed[31:0]    reg_psum_34_15;
wire signed[31:0]    reg_weight_34_16;
wire signed[31:0]    reg_psum_34_16;
wire signed[31:0]    reg_weight_34_17;
wire signed[31:0]    reg_psum_34_17;
wire signed[31:0]    reg_weight_34_18;
wire signed[31:0]    reg_psum_34_18;
wire signed[31:0]    reg_weight_34_19;
wire signed[31:0]    reg_psum_34_19;
wire signed[31:0]    reg_weight_34_20;
wire signed[31:0]    reg_psum_34_20;
wire signed[31:0]    reg_weight_34_21;
wire signed[31:0]    reg_psum_34_21;
wire signed[31:0]    reg_weight_34_22;
wire signed[31:0]    reg_psum_34_22;
wire signed[31:0]    reg_weight_34_23;
wire signed[31:0]    reg_psum_34_23;
wire signed[31:0]    reg_weight_34_24;
wire signed[31:0]    reg_psum_34_24;
wire signed[31:0]    reg_weight_34_25;
wire signed[31:0]    reg_psum_34_25;
wire signed[31:0]    reg_weight_34_26;
wire signed[31:0]    reg_psum_34_26;
wire signed[31:0]    reg_weight_34_27;
wire signed[31:0]    reg_psum_34_27;
wire signed[31:0]    reg_weight_34_28;
wire signed[31:0]    reg_psum_34_28;
wire signed[31:0]    reg_weight_34_29;
wire signed[31:0]    reg_psum_34_29;
wire signed[31:0]    reg_weight_34_30;
wire signed[31:0]    reg_psum_34_30;
wire signed[31:0]    reg_weight_34_31;
wire signed[31:0]    reg_psum_34_31;
wire signed[31:0]    reg_weight_34_32;
wire signed[31:0]    reg_psum_34_32;
wire signed[31:0]    reg_weight_34_33;
wire signed[31:0]    reg_psum_34_33;
wire signed[31:0]    reg_weight_34_34;
wire signed[31:0]    reg_psum_34_34;
wire signed[31:0]    reg_weight_34_35;
wire signed[31:0]    reg_psum_34_35;
wire signed[31:0]    reg_weight_34_36;
wire signed[31:0]    reg_psum_34_36;
wire signed[31:0]    reg_weight_34_37;
wire signed[31:0]    reg_psum_34_37;
wire signed[31:0]    reg_weight_34_38;
wire signed[31:0]    reg_psum_34_38;
wire signed[31:0]    reg_weight_34_39;
wire signed[31:0]    reg_psum_34_39;
wire signed[31:0]    reg_weight_34_40;
wire signed[31:0]    reg_psum_34_40;
wire signed[31:0]    reg_weight_34_41;
wire signed[31:0]    reg_psum_34_41;
wire signed[31:0]    reg_weight_34_42;
wire signed[31:0]    reg_psum_34_42;
wire signed[31:0]    reg_weight_34_43;
wire signed[31:0]    reg_psum_34_43;
wire signed[31:0]    reg_weight_34_44;
wire signed[31:0]    reg_psum_34_44;
wire signed[31:0]    reg_weight_34_45;
wire signed[31:0]    reg_psum_34_45;
wire signed[31:0]    reg_weight_34_46;
wire signed[31:0]    reg_psum_34_46;
wire signed[31:0]    reg_weight_34_47;
wire signed[31:0]    reg_psum_34_47;
wire signed[31:0]    reg_weight_34_48;
wire signed[31:0]    reg_psum_34_48;
wire signed[31:0]    reg_weight_34_49;
wire signed[31:0]    reg_psum_34_49;
wire signed[31:0]    reg_weight_34_50;
wire signed[31:0]    reg_psum_34_50;
wire signed[31:0]    reg_weight_34_51;
wire signed[31:0]    reg_psum_34_51;
wire signed[31:0]    reg_weight_34_52;
wire signed[31:0]    reg_psum_34_52;
wire signed[31:0]    reg_weight_34_53;
wire signed[31:0]    reg_psum_34_53;
wire signed[31:0]    reg_weight_34_54;
wire signed[31:0]    reg_psum_34_54;
wire signed[31:0]    reg_weight_34_55;
wire signed[31:0]    reg_psum_34_55;
wire signed[31:0]    reg_weight_34_56;
wire signed[31:0]    reg_psum_34_56;
wire signed[31:0]    reg_weight_34_57;
wire signed[31:0]    reg_psum_34_57;
wire signed[31:0]    reg_weight_34_58;
wire signed[31:0]    reg_psum_34_58;
wire signed[31:0]    reg_weight_34_59;
wire signed[31:0]    reg_psum_34_59;
wire signed[31:0]    reg_weight_34_60;
wire signed[31:0]    reg_psum_34_60;
wire signed[31:0]    reg_weight_34_61;
wire signed[31:0]    reg_psum_34_61;
wire signed[31:0]    reg_weight_34_62;
wire signed[31:0]    reg_psum_34_62;
wire signed[31:0]    reg_weight_34_63;
wire signed[31:0]    reg_psum_34_63;
wire signed[31:0]    reg_weight_35_0;
wire signed[31:0]    reg_psum_35_0;
wire signed[31:0]    reg_weight_35_1;
wire signed[31:0]    reg_psum_35_1;
wire signed[31:0]    reg_weight_35_2;
wire signed[31:0]    reg_psum_35_2;
wire signed[31:0]    reg_weight_35_3;
wire signed[31:0]    reg_psum_35_3;
wire signed[31:0]    reg_weight_35_4;
wire signed[31:0]    reg_psum_35_4;
wire signed[31:0]    reg_weight_35_5;
wire signed[31:0]    reg_psum_35_5;
wire signed[31:0]    reg_weight_35_6;
wire signed[31:0]    reg_psum_35_6;
wire signed[31:0]    reg_weight_35_7;
wire signed[31:0]    reg_psum_35_7;
wire signed[31:0]    reg_weight_35_8;
wire signed[31:0]    reg_psum_35_8;
wire signed[31:0]    reg_weight_35_9;
wire signed[31:0]    reg_psum_35_9;
wire signed[31:0]    reg_weight_35_10;
wire signed[31:0]    reg_psum_35_10;
wire signed[31:0]    reg_weight_35_11;
wire signed[31:0]    reg_psum_35_11;
wire signed[31:0]    reg_weight_35_12;
wire signed[31:0]    reg_psum_35_12;
wire signed[31:0]    reg_weight_35_13;
wire signed[31:0]    reg_psum_35_13;
wire signed[31:0]    reg_weight_35_14;
wire signed[31:0]    reg_psum_35_14;
wire signed[31:0]    reg_weight_35_15;
wire signed[31:0]    reg_psum_35_15;
wire signed[31:0]    reg_weight_35_16;
wire signed[31:0]    reg_psum_35_16;
wire signed[31:0]    reg_weight_35_17;
wire signed[31:0]    reg_psum_35_17;
wire signed[31:0]    reg_weight_35_18;
wire signed[31:0]    reg_psum_35_18;
wire signed[31:0]    reg_weight_35_19;
wire signed[31:0]    reg_psum_35_19;
wire signed[31:0]    reg_weight_35_20;
wire signed[31:0]    reg_psum_35_20;
wire signed[31:0]    reg_weight_35_21;
wire signed[31:0]    reg_psum_35_21;
wire signed[31:0]    reg_weight_35_22;
wire signed[31:0]    reg_psum_35_22;
wire signed[31:0]    reg_weight_35_23;
wire signed[31:0]    reg_psum_35_23;
wire signed[31:0]    reg_weight_35_24;
wire signed[31:0]    reg_psum_35_24;
wire signed[31:0]    reg_weight_35_25;
wire signed[31:0]    reg_psum_35_25;
wire signed[31:0]    reg_weight_35_26;
wire signed[31:0]    reg_psum_35_26;
wire signed[31:0]    reg_weight_35_27;
wire signed[31:0]    reg_psum_35_27;
wire signed[31:0]    reg_weight_35_28;
wire signed[31:0]    reg_psum_35_28;
wire signed[31:0]    reg_weight_35_29;
wire signed[31:0]    reg_psum_35_29;
wire signed[31:0]    reg_weight_35_30;
wire signed[31:0]    reg_psum_35_30;
wire signed[31:0]    reg_weight_35_31;
wire signed[31:0]    reg_psum_35_31;
wire signed[31:0]    reg_weight_35_32;
wire signed[31:0]    reg_psum_35_32;
wire signed[31:0]    reg_weight_35_33;
wire signed[31:0]    reg_psum_35_33;
wire signed[31:0]    reg_weight_35_34;
wire signed[31:0]    reg_psum_35_34;
wire signed[31:0]    reg_weight_35_35;
wire signed[31:0]    reg_psum_35_35;
wire signed[31:0]    reg_weight_35_36;
wire signed[31:0]    reg_psum_35_36;
wire signed[31:0]    reg_weight_35_37;
wire signed[31:0]    reg_psum_35_37;
wire signed[31:0]    reg_weight_35_38;
wire signed[31:0]    reg_psum_35_38;
wire signed[31:0]    reg_weight_35_39;
wire signed[31:0]    reg_psum_35_39;
wire signed[31:0]    reg_weight_35_40;
wire signed[31:0]    reg_psum_35_40;
wire signed[31:0]    reg_weight_35_41;
wire signed[31:0]    reg_psum_35_41;
wire signed[31:0]    reg_weight_35_42;
wire signed[31:0]    reg_psum_35_42;
wire signed[31:0]    reg_weight_35_43;
wire signed[31:0]    reg_psum_35_43;
wire signed[31:0]    reg_weight_35_44;
wire signed[31:0]    reg_psum_35_44;
wire signed[31:0]    reg_weight_35_45;
wire signed[31:0]    reg_psum_35_45;
wire signed[31:0]    reg_weight_35_46;
wire signed[31:0]    reg_psum_35_46;
wire signed[31:0]    reg_weight_35_47;
wire signed[31:0]    reg_psum_35_47;
wire signed[31:0]    reg_weight_35_48;
wire signed[31:0]    reg_psum_35_48;
wire signed[31:0]    reg_weight_35_49;
wire signed[31:0]    reg_psum_35_49;
wire signed[31:0]    reg_weight_35_50;
wire signed[31:0]    reg_psum_35_50;
wire signed[31:0]    reg_weight_35_51;
wire signed[31:0]    reg_psum_35_51;
wire signed[31:0]    reg_weight_35_52;
wire signed[31:0]    reg_psum_35_52;
wire signed[31:0]    reg_weight_35_53;
wire signed[31:0]    reg_psum_35_53;
wire signed[31:0]    reg_weight_35_54;
wire signed[31:0]    reg_psum_35_54;
wire signed[31:0]    reg_weight_35_55;
wire signed[31:0]    reg_psum_35_55;
wire signed[31:0]    reg_weight_35_56;
wire signed[31:0]    reg_psum_35_56;
wire signed[31:0]    reg_weight_35_57;
wire signed[31:0]    reg_psum_35_57;
wire signed[31:0]    reg_weight_35_58;
wire signed[31:0]    reg_psum_35_58;
wire signed[31:0]    reg_weight_35_59;
wire signed[31:0]    reg_psum_35_59;
wire signed[31:0]    reg_weight_35_60;
wire signed[31:0]    reg_psum_35_60;
wire signed[31:0]    reg_weight_35_61;
wire signed[31:0]    reg_psum_35_61;
wire signed[31:0]    reg_weight_35_62;
wire signed[31:0]    reg_psum_35_62;
wire signed[31:0]    reg_weight_35_63;
wire signed[31:0]    reg_psum_35_63;
wire signed[31:0]    reg_weight_36_0;
wire signed[31:0]    reg_psum_36_0;
wire signed[31:0]    reg_weight_36_1;
wire signed[31:0]    reg_psum_36_1;
wire signed[31:0]    reg_weight_36_2;
wire signed[31:0]    reg_psum_36_2;
wire signed[31:0]    reg_weight_36_3;
wire signed[31:0]    reg_psum_36_3;
wire signed[31:0]    reg_weight_36_4;
wire signed[31:0]    reg_psum_36_4;
wire signed[31:0]    reg_weight_36_5;
wire signed[31:0]    reg_psum_36_5;
wire signed[31:0]    reg_weight_36_6;
wire signed[31:0]    reg_psum_36_6;
wire signed[31:0]    reg_weight_36_7;
wire signed[31:0]    reg_psum_36_7;
wire signed[31:0]    reg_weight_36_8;
wire signed[31:0]    reg_psum_36_8;
wire signed[31:0]    reg_weight_36_9;
wire signed[31:0]    reg_psum_36_9;
wire signed[31:0]    reg_weight_36_10;
wire signed[31:0]    reg_psum_36_10;
wire signed[31:0]    reg_weight_36_11;
wire signed[31:0]    reg_psum_36_11;
wire signed[31:0]    reg_weight_36_12;
wire signed[31:0]    reg_psum_36_12;
wire signed[31:0]    reg_weight_36_13;
wire signed[31:0]    reg_psum_36_13;
wire signed[31:0]    reg_weight_36_14;
wire signed[31:0]    reg_psum_36_14;
wire signed[31:0]    reg_weight_36_15;
wire signed[31:0]    reg_psum_36_15;
wire signed[31:0]    reg_weight_36_16;
wire signed[31:0]    reg_psum_36_16;
wire signed[31:0]    reg_weight_36_17;
wire signed[31:0]    reg_psum_36_17;
wire signed[31:0]    reg_weight_36_18;
wire signed[31:0]    reg_psum_36_18;
wire signed[31:0]    reg_weight_36_19;
wire signed[31:0]    reg_psum_36_19;
wire signed[31:0]    reg_weight_36_20;
wire signed[31:0]    reg_psum_36_20;
wire signed[31:0]    reg_weight_36_21;
wire signed[31:0]    reg_psum_36_21;
wire signed[31:0]    reg_weight_36_22;
wire signed[31:0]    reg_psum_36_22;
wire signed[31:0]    reg_weight_36_23;
wire signed[31:0]    reg_psum_36_23;
wire signed[31:0]    reg_weight_36_24;
wire signed[31:0]    reg_psum_36_24;
wire signed[31:0]    reg_weight_36_25;
wire signed[31:0]    reg_psum_36_25;
wire signed[31:0]    reg_weight_36_26;
wire signed[31:0]    reg_psum_36_26;
wire signed[31:0]    reg_weight_36_27;
wire signed[31:0]    reg_psum_36_27;
wire signed[31:0]    reg_weight_36_28;
wire signed[31:0]    reg_psum_36_28;
wire signed[31:0]    reg_weight_36_29;
wire signed[31:0]    reg_psum_36_29;
wire signed[31:0]    reg_weight_36_30;
wire signed[31:0]    reg_psum_36_30;
wire signed[31:0]    reg_weight_36_31;
wire signed[31:0]    reg_psum_36_31;
wire signed[31:0]    reg_weight_36_32;
wire signed[31:0]    reg_psum_36_32;
wire signed[31:0]    reg_weight_36_33;
wire signed[31:0]    reg_psum_36_33;
wire signed[31:0]    reg_weight_36_34;
wire signed[31:0]    reg_psum_36_34;
wire signed[31:0]    reg_weight_36_35;
wire signed[31:0]    reg_psum_36_35;
wire signed[31:0]    reg_weight_36_36;
wire signed[31:0]    reg_psum_36_36;
wire signed[31:0]    reg_weight_36_37;
wire signed[31:0]    reg_psum_36_37;
wire signed[31:0]    reg_weight_36_38;
wire signed[31:0]    reg_psum_36_38;
wire signed[31:0]    reg_weight_36_39;
wire signed[31:0]    reg_psum_36_39;
wire signed[31:0]    reg_weight_36_40;
wire signed[31:0]    reg_psum_36_40;
wire signed[31:0]    reg_weight_36_41;
wire signed[31:0]    reg_psum_36_41;
wire signed[31:0]    reg_weight_36_42;
wire signed[31:0]    reg_psum_36_42;
wire signed[31:0]    reg_weight_36_43;
wire signed[31:0]    reg_psum_36_43;
wire signed[31:0]    reg_weight_36_44;
wire signed[31:0]    reg_psum_36_44;
wire signed[31:0]    reg_weight_36_45;
wire signed[31:0]    reg_psum_36_45;
wire signed[31:0]    reg_weight_36_46;
wire signed[31:0]    reg_psum_36_46;
wire signed[31:0]    reg_weight_36_47;
wire signed[31:0]    reg_psum_36_47;
wire signed[31:0]    reg_weight_36_48;
wire signed[31:0]    reg_psum_36_48;
wire signed[31:0]    reg_weight_36_49;
wire signed[31:0]    reg_psum_36_49;
wire signed[31:0]    reg_weight_36_50;
wire signed[31:0]    reg_psum_36_50;
wire signed[31:0]    reg_weight_36_51;
wire signed[31:0]    reg_psum_36_51;
wire signed[31:0]    reg_weight_36_52;
wire signed[31:0]    reg_psum_36_52;
wire signed[31:0]    reg_weight_36_53;
wire signed[31:0]    reg_psum_36_53;
wire signed[31:0]    reg_weight_36_54;
wire signed[31:0]    reg_psum_36_54;
wire signed[31:0]    reg_weight_36_55;
wire signed[31:0]    reg_psum_36_55;
wire signed[31:0]    reg_weight_36_56;
wire signed[31:0]    reg_psum_36_56;
wire signed[31:0]    reg_weight_36_57;
wire signed[31:0]    reg_psum_36_57;
wire signed[31:0]    reg_weight_36_58;
wire signed[31:0]    reg_psum_36_58;
wire signed[31:0]    reg_weight_36_59;
wire signed[31:0]    reg_psum_36_59;
wire signed[31:0]    reg_weight_36_60;
wire signed[31:0]    reg_psum_36_60;
wire signed[31:0]    reg_weight_36_61;
wire signed[31:0]    reg_psum_36_61;
wire signed[31:0]    reg_weight_36_62;
wire signed[31:0]    reg_psum_36_62;
wire signed[31:0]    reg_weight_36_63;
wire signed[31:0]    reg_psum_36_63;
wire signed[31:0]    reg_weight_37_0;
wire signed[31:0]    reg_psum_37_0;
wire signed[31:0]    reg_weight_37_1;
wire signed[31:0]    reg_psum_37_1;
wire signed[31:0]    reg_weight_37_2;
wire signed[31:0]    reg_psum_37_2;
wire signed[31:0]    reg_weight_37_3;
wire signed[31:0]    reg_psum_37_3;
wire signed[31:0]    reg_weight_37_4;
wire signed[31:0]    reg_psum_37_4;
wire signed[31:0]    reg_weight_37_5;
wire signed[31:0]    reg_psum_37_5;
wire signed[31:0]    reg_weight_37_6;
wire signed[31:0]    reg_psum_37_6;
wire signed[31:0]    reg_weight_37_7;
wire signed[31:0]    reg_psum_37_7;
wire signed[31:0]    reg_weight_37_8;
wire signed[31:0]    reg_psum_37_8;
wire signed[31:0]    reg_weight_37_9;
wire signed[31:0]    reg_psum_37_9;
wire signed[31:0]    reg_weight_37_10;
wire signed[31:0]    reg_psum_37_10;
wire signed[31:0]    reg_weight_37_11;
wire signed[31:0]    reg_psum_37_11;
wire signed[31:0]    reg_weight_37_12;
wire signed[31:0]    reg_psum_37_12;
wire signed[31:0]    reg_weight_37_13;
wire signed[31:0]    reg_psum_37_13;
wire signed[31:0]    reg_weight_37_14;
wire signed[31:0]    reg_psum_37_14;
wire signed[31:0]    reg_weight_37_15;
wire signed[31:0]    reg_psum_37_15;
wire signed[31:0]    reg_weight_37_16;
wire signed[31:0]    reg_psum_37_16;
wire signed[31:0]    reg_weight_37_17;
wire signed[31:0]    reg_psum_37_17;
wire signed[31:0]    reg_weight_37_18;
wire signed[31:0]    reg_psum_37_18;
wire signed[31:0]    reg_weight_37_19;
wire signed[31:0]    reg_psum_37_19;
wire signed[31:0]    reg_weight_37_20;
wire signed[31:0]    reg_psum_37_20;
wire signed[31:0]    reg_weight_37_21;
wire signed[31:0]    reg_psum_37_21;
wire signed[31:0]    reg_weight_37_22;
wire signed[31:0]    reg_psum_37_22;
wire signed[31:0]    reg_weight_37_23;
wire signed[31:0]    reg_psum_37_23;
wire signed[31:0]    reg_weight_37_24;
wire signed[31:0]    reg_psum_37_24;
wire signed[31:0]    reg_weight_37_25;
wire signed[31:0]    reg_psum_37_25;
wire signed[31:0]    reg_weight_37_26;
wire signed[31:0]    reg_psum_37_26;
wire signed[31:0]    reg_weight_37_27;
wire signed[31:0]    reg_psum_37_27;
wire signed[31:0]    reg_weight_37_28;
wire signed[31:0]    reg_psum_37_28;
wire signed[31:0]    reg_weight_37_29;
wire signed[31:0]    reg_psum_37_29;
wire signed[31:0]    reg_weight_37_30;
wire signed[31:0]    reg_psum_37_30;
wire signed[31:0]    reg_weight_37_31;
wire signed[31:0]    reg_psum_37_31;
wire signed[31:0]    reg_weight_37_32;
wire signed[31:0]    reg_psum_37_32;
wire signed[31:0]    reg_weight_37_33;
wire signed[31:0]    reg_psum_37_33;
wire signed[31:0]    reg_weight_37_34;
wire signed[31:0]    reg_psum_37_34;
wire signed[31:0]    reg_weight_37_35;
wire signed[31:0]    reg_psum_37_35;
wire signed[31:0]    reg_weight_37_36;
wire signed[31:0]    reg_psum_37_36;
wire signed[31:0]    reg_weight_37_37;
wire signed[31:0]    reg_psum_37_37;
wire signed[31:0]    reg_weight_37_38;
wire signed[31:0]    reg_psum_37_38;
wire signed[31:0]    reg_weight_37_39;
wire signed[31:0]    reg_psum_37_39;
wire signed[31:0]    reg_weight_37_40;
wire signed[31:0]    reg_psum_37_40;
wire signed[31:0]    reg_weight_37_41;
wire signed[31:0]    reg_psum_37_41;
wire signed[31:0]    reg_weight_37_42;
wire signed[31:0]    reg_psum_37_42;
wire signed[31:0]    reg_weight_37_43;
wire signed[31:0]    reg_psum_37_43;
wire signed[31:0]    reg_weight_37_44;
wire signed[31:0]    reg_psum_37_44;
wire signed[31:0]    reg_weight_37_45;
wire signed[31:0]    reg_psum_37_45;
wire signed[31:0]    reg_weight_37_46;
wire signed[31:0]    reg_psum_37_46;
wire signed[31:0]    reg_weight_37_47;
wire signed[31:0]    reg_psum_37_47;
wire signed[31:0]    reg_weight_37_48;
wire signed[31:0]    reg_psum_37_48;
wire signed[31:0]    reg_weight_37_49;
wire signed[31:0]    reg_psum_37_49;
wire signed[31:0]    reg_weight_37_50;
wire signed[31:0]    reg_psum_37_50;
wire signed[31:0]    reg_weight_37_51;
wire signed[31:0]    reg_psum_37_51;
wire signed[31:0]    reg_weight_37_52;
wire signed[31:0]    reg_psum_37_52;
wire signed[31:0]    reg_weight_37_53;
wire signed[31:0]    reg_psum_37_53;
wire signed[31:0]    reg_weight_37_54;
wire signed[31:0]    reg_psum_37_54;
wire signed[31:0]    reg_weight_37_55;
wire signed[31:0]    reg_psum_37_55;
wire signed[31:0]    reg_weight_37_56;
wire signed[31:0]    reg_psum_37_56;
wire signed[31:0]    reg_weight_37_57;
wire signed[31:0]    reg_psum_37_57;
wire signed[31:0]    reg_weight_37_58;
wire signed[31:0]    reg_psum_37_58;
wire signed[31:0]    reg_weight_37_59;
wire signed[31:0]    reg_psum_37_59;
wire signed[31:0]    reg_weight_37_60;
wire signed[31:0]    reg_psum_37_60;
wire signed[31:0]    reg_weight_37_61;
wire signed[31:0]    reg_psum_37_61;
wire signed[31:0]    reg_weight_37_62;
wire signed[31:0]    reg_psum_37_62;
wire signed[31:0]    reg_weight_37_63;
wire signed[31:0]    reg_psum_37_63;
wire signed[31:0]    reg_weight_38_0;
wire signed[31:0]    reg_psum_38_0;
wire signed[31:0]    reg_weight_38_1;
wire signed[31:0]    reg_psum_38_1;
wire signed[31:0]    reg_weight_38_2;
wire signed[31:0]    reg_psum_38_2;
wire signed[31:0]    reg_weight_38_3;
wire signed[31:0]    reg_psum_38_3;
wire signed[31:0]    reg_weight_38_4;
wire signed[31:0]    reg_psum_38_4;
wire signed[31:0]    reg_weight_38_5;
wire signed[31:0]    reg_psum_38_5;
wire signed[31:0]    reg_weight_38_6;
wire signed[31:0]    reg_psum_38_6;
wire signed[31:0]    reg_weight_38_7;
wire signed[31:0]    reg_psum_38_7;
wire signed[31:0]    reg_weight_38_8;
wire signed[31:0]    reg_psum_38_8;
wire signed[31:0]    reg_weight_38_9;
wire signed[31:0]    reg_psum_38_9;
wire signed[31:0]    reg_weight_38_10;
wire signed[31:0]    reg_psum_38_10;
wire signed[31:0]    reg_weight_38_11;
wire signed[31:0]    reg_psum_38_11;
wire signed[31:0]    reg_weight_38_12;
wire signed[31:0]    reg_psum_38_12;
wire signed[31:0]    reg_weight_38_13;
wire signed[31:0]    reg_psum_38_13;
wire signed[31:0]    reg_weight_38_14;
wire signed[31:0]    reg_psum_38_14;
wire signed[31:0]    reg_weight_38_15;
wire signed[31:0]    reg_psum_38_15;
wire signed[31:0]    reg_weight_38_16;
wire signed[31:0]    reg_psum_38_16;
wire signed[31:0]    reg_weight_38_17;
wire signed[31:0]    reg_psum_38_17;
wire signed[31:0]    reg_weight_38_18;
wire signed[31:0]    reg_psum_38_18;
wire signed[31:0]    reg_weight_38_19;
wire signed[31:0]    reg_psum_38_19;
wire signed[31:0]    reg_weight_38_20;
wire signed[31:0]    reg_psum_38_20;
wire signed[31:0]    reg_weight_38_21;
wire signed[31:0]    reg_psum_38_21;
wire signed[31:0]    reg_weight_38_22;
wire signed[31:0]    reg_psum_38_22;
wire signed[31:0]    reg_weight_38_23;
wire signed[31:0]    reg_psum_38_23;
wire signed[31:0]    reg_weight_38_24;
wire signed[31:0]    reg_psum_38_24;
wire signed[31:0]    reg_weight_38_25;
wire signed[31:0]    reg_psum_38_25;
wire signed[31:0]    reg_weight_38_26;
wire signed[31:0]    reg_psum_38_26;
wire signed[31:0]    reg_weight_38_27;
wire signed[31:0]    reg_psum_38_27;
wire signed[31:0]    reg_weight_38_28;
wire signed[31:0]    reg_psum_38_28;
wire signed[31:0]    reg_weight_38_29;
wire signed[31:0]    reg_psum_38_29;
wire signed[31:0]    reg_weight_38_30;
wire signed[31:0]    reg_psum_38_30;
wire signed[31:0]    reg_weight_38_31;
wire signed[31:0]    reg_psum_38_31;
wire signed[31:0]    reg_weight_38_32;
wire signed[31:0]    reg_psum_38_32;
wire signed[31:0]    reg_weight_38_33;
wire signed[31:0]    reg_psum_38_33;
wire signed[31:0]    reg_weight_38_34;
wire signed[31:0]    reg_psum_38_34;
wire signed[31:0]    reg_weight_38_35;
wire signed[31:0]    reg_psum_38_35;
wire signed[31:0]    reg_weight_38_36;
wire signed[31:0]    reg_psum_38_36;
wire signed[31:0]    reg_weight_38_37;
wire signed[31:0]    reg_psum_38_37;
wire signed[31:0]    reg_weight_38_38;
wire signed[31:0]    reg_psum_38_38;
wire signed[31:0]    reg_weight_38_39;
wire signed[31:0]    reg_psum_38_39;
wire signed[31:0]    reg_weight_38_40;
wire signed[31:0]    reg_psum_38_40;
wire signed[31:0]    reg_weight_38_41;
wire signed[31:0]    reg_psum_38_41;
wire signed[31:0]    reg_weight_38_42;
wire signed[31:0]    reg_psum_38_42;
wire signed[31:0]    reg_weight_38_43;
wire signed[31:0]    reg_psum_38_43;
wire signed[31:0]    reg_weight_38_44;
wire signed[31:0]    reg_psum_38_44;
wire signed[31:0]    reg_weight_38_45;
wire signed[31:0]    reg_psum_38_45;
wire signed[31:0]    reg_weight_38_46;
wire signed[31:0]    reg_psum_38_46;
wire signed[31:0]    reg_weight_38_47;
wire signed[31:0]    reg_psum_38_47;
wire signed[31:0]    reg_weight_38_48;
wire signed[31:0]    reg_psum_38_48;
wire signed[31:0]    reg_weight_38_49;
wire signed[31:0]    reg_psum_38_49;
wire signed[31:0]    reg_weight_38_50;
wire signed[31:0]    reg_psum_38_50;
wire signed[31:0]    reg_weight_38_51;
wire signed[31:0]    reg_psum_38_51;
wire signed[31:0]    reg_weight_38_52;
wire signed[31:0]    reg_psum_38_52;
wire signed[31:0]    reg_weight_38_53;
wire signed[31:0]    reg_psum_38_53;
wire signed[31:0]    reg_weight_38_54;
wire signed[31:0]    reg_psum_38_54;
wire signed[31:0]    reg_weight_38_55;
wire signed[31:0]    reg_psum_38_55;
wire signed[31:0]    reg_weight_38_56;
wire signed[31:0]    reg_psum_38_56;
wire signed[31:0]    reg_weight_38_57;
wire signed[31:0]    reg_psum_38_57;
wire signed[31:0]    reg_weight_38_58;
wire signed[31:0]    reg_psum_38_58;
wire signed[31:0]    reg_weight_38_59;
wire signed[31:0]    reg_psum_38_59;
wire signed[31:0]    reg_weight_38_60;
wire signed[31:0]    reg_psum_38_60;
wire signed[31:0]    reg_weight_38_61;
wire signed[31:0]    reg_psum_38_61;
wire signed[31:0]    reg_weight_38_62;
wire signed[31:0]    reg_psum_38_62;
wire signed[31:0]    reg_weight_38_63;
wire signed[31:0]    reg_psum_38_63;
wire signed[31:0]    reg_weight_39_0;
wire signed[31:0]    reg_psum_39_0;
wire signed[31:0]    reg_weight_39_1;
wire signed[31:0]    reg_psum_39_1;
wire signed[31:0]    reg_weight_39_2;
wire signed[31:0]    reg_psum_39_2;
wire signed[31:0]    reg_weight_39_3;
wire signed[31:0]    reg_psum_39_3;
wire signed[31:0]    reg_weight_39_4;
wire signed[31:0]    reg_psum_39_4;
wire signed[31:0]    reg_weight_39_5;
wire signed[31:0]    reg_psum_39_5;
wire signed[31:0]    reg_weight_39_6;
wire signed[31:0]    reg_psum_39_6;
wire signed[31:0]    reg_weight_39_7;
wire signed[31:0]    reg_psum_39_7;
wire signed[31:0]    reg_weight_39_8;
wire signed[31:0]    reg_psum_39_8;
wire signed[31:0]    reg_weight_39_9;
wire signed[31:0]    reg_psum_39_9;
wire signed[31:0]    reg_weight_39_10;
wire signed[31:0]    reg_psum_39_10;
wire signed[31:0]    reg_weight_39_11;
wire signed[31:0]    reg_psum_39_11;
wire signed[31:0]    reg_weight_39_12;
wire signed[31:0]    reg_psum_39_12;
wire signed[31:0]    reg_weight_39_13;
wire signed[31:0]    reg_psum_39_13;
wire signed[31:0]    reg_weight_39_14;
wire signed[31:0]    reg_psum_39_14;
wire signed[31:0]    reg_weight_39_15;
wire signed[31:0]    reg_psum_39_15;
wire signed[31:0]    reg_weight_39_16;
wire signed[31:0]    reg_psum_39_16;
wire signed[31:0]    reg_weight_39_17;
wire signed[31:0]    reg_psum_39_17;
wire signed[31:0]    reg_weight_39_18;
wire signed[31:0]    reg_psum_39_18;
wire signed[31:0]    reg_weight_39_19;
wire signed[31:0]    reg_psum_39_19;
wire signed[31:0]    reg_weight_39_20;
wire signed[31:0]    reg_psum_39_20;
wire signed[31:0]    reg_weight_39_21;
wire signed[31:0]    reg_psum_39_21;
wire signed[31:0]    reg_weight_39_22;
wire signed[31:0]    reg_psum_39_22;
wire signed[31:0]    reg_weight_39_23;
wire signed[31:0]    reg_psum_39_23;
wire signed[31:0]    reg_weight_39_24;
wire signed[31:0]    reg_psum_39_24;
wire signed[31:0]    reg_weight_39_25;
wire signed[31:0]    reg_psum_39_25;
wire signed[31:0]    reg_weight_39_26;
wire signed[31:0]    reg_psum_39_26;
wire signed[31:0]    reg_weight_39_27;
wire signed[31:0]    reg_psum_39_27;
wire signed[31:0]    reg_weight_39_28;
wire signed[31:0]    reg_psum_39_28;
wire signed[31:0]    reg_weight_39_29;
wire signed[31:0]    reg_psum_39_29;
wire signed[31:0]    reg_weight_39_30;
wire signed[31:0]    reg_psum_39_30;
wire signed[31:0]    reg_weight_39_31;
wire signed[31:0]    reg_psum_39_31;
wire signed[31:0]    reg_weight_39_32;
wire signed[31:0]    reg_psum_39_32;
wire signed[31:0]    reg_weight_39_33;
wire signed[31:0]    reg_psum_39_33;
wire signed[31:0]    reg_weight_39_34;
wire signed[31:0]    reg_psum_39_34;
wire signed[31:0]    reg_weight_39_35;
wire signed[31:0]    reg_psum_39_35;
wire signed[31:0]    reg_weight_39_36;
wire signed[31:0]    reg_psum_39_36;
wire signed[31:0]    reg_weight_39_37;
wire signed[31:0]    reg_psum_39_37;
wire signed[31:0]    reg_weight_39_38;
wire signed[31:0]    reg_psum_39_38;
wire signed[31:0]    reg_weight_39_39;
wire signed[31:0]    reg_psum_39_39;
wire signed[31:0]    reg_weight_39_40;
wire signed[31:0]    reg_psum_39_40;
wire signed[31:0]    reg_weight_39_41;
wire signed[31:0]    reg_psum_39_41;
wire signed[31:0]    reg_weight_39_42;
wire signed[31:0]    reg_psum_39_42;
wire signed[31:0]    reg_weight_39_43;
wire signed[31:0]    reg_psum_39_43;
wire signed[31:0]    reg_weight_39_44;
wire signed[31:0]    reg_psum_39_44;
wire signed[31:0]    reg_weight_39_45;
wire signed[31:0]    reg_psum_39_45;
wire signed[31:0]    reg_weight_39_46;
wire signed[31:0]    reg_psum_39_46;
wire signed[31:0]    reg_weight_39_47;
wire signed[31:0]    reg_psum_39_47;
wire signed[31:0]    reg_weight_39_48;
wire signed[31:0]    reg_psum_39_48;
wire signed[31:0]    reg_weight_39_49;
wire signed[31:0]    reg_psum_39_49;
wire signed[31:0]    reg_weight_39_50;
wire signed[31:0]    reg_psum_39_50;
wire signed[31:0]    reg_weight_39_51;
wire signed[31:0]    reg_psum_39_51;
wire signed[31:0]    reg_weight_39_52;
wire signed[31:0]    reg_psum_39_52;
wire signed[31:0]    reg_weight_39_53;
wire signed[31:0]    reg_psum_39_53;
wire signed[31:0]    reg_weight_39_54;
wire signed[31:0]    reg_psum_39_54;
wire signed[31:0]    reg_weight_39_55;
wire signed[31:0]    reg_psum_39_55;
wire signed[31:0]    reg_weight_39_56;
wire signed[31:0]    reg_psum_39_56;
wire signed[31:0]    reg_weight_39_57;
wire signed[31:0]    reg_psum_39_57;
wire signed[31:0]    reg_weight_39_58;
wire signed[31:0]    reg_psum_39_58;
wire signed[31:0]    reg_weight_39_59;
wire signed[31:0]    reg_psum_39_59;
wire signed[31:0]    reg_weight_39_60;
wire signed[31:0]    reg_psum_39_60;
wire signed[31:0]    reg_weight_39_61;
wire signed[31:0]    reg_psum_39_61;
wire signed[31:0]    reg_weight_39_62;
wire signed[31:0]    reg_psum_39_62;
wire signed[31:0]    reg_weight_39_63;
wire signed[31:0]    reg_psum_39_63;
wire signed[31:0]    reg_weight_40_0;
wire signed[31:0]    reg_psum_40_0;
wire signed[31:0]    reg_weight_40_1;
wire signed[31:0]    reg_psum_40_1;
wire signed[31:0]    reg_weight_40_2;
wire signed[31:0]    reg_psum_40_2;
wire signed[31:0]    reg_weight_40_3;
wire signed[31:0]    reg_psum_40_3;
wire signed[31:0]    reg_weight_40_4;
wire signed[31:0]    reg_psum_40_4;
wire signed[31:0]    reg_weight_40_5;
wire signed[31:0]    reg_psum_40_5;
wire signed[31:0]    reg_weight_40_6;
wire signed[31:0]    reg_psum_40_6;
wire signed[31:0]    reg_weight_40_7;
wire signed[31:0]    reg_psum_40_7;
wire signed[31:0]    reg_weight_40_8;
wire signed[31:0]    reg_psum_40_8;
wire signed[31:0]    reg_weight_40_9;
wire signed[31:0]    reg_psum_40_9;
wire signed[31:0]    reg_weight_40_10;
wire signed[31:0]    reg_psum_40_10;
wire signed[31:0]    reg_weight_40_11;
wire signed[31:0]    reg_psum_40_11;
wire signed[31:0]    reg_weight_40_12;
wire signed[31:0]    reg_psum_40_12;
wire signed[31:0]    reg_weight_40_13;
wire signed[31:0]    reg_psum_40_13;
wire signed[31:0]    reg_weight_40_14;
wire signed[31:0]    reg_psum_40_14;
wire signed[31:0]    reg_weight_40_15;
wire signed[31:0]    reg_psum_40_15;
wire signed[31:0]    reg_weight_40_16;
wire signed[31:0]    reg_psum_40_16;
wire signed[31:0]    reg_weight_40_17;
wire signed[31:0]    reg_psum_40_17;
wire signed[31:0]    reg_weight_40_18;
wire signed[31:0]    reg_psum_40_18;
wire signed[31:0]    reg_weight_40_19;
wire signed[31:0]    reg_psum_40_19;
wire signed[31:0]    reg_weight_40_20;
wire signed[31:0]    reg_psum_40_20;
wire signed[31:0]    reg_weight_40_21;
wire signed[31:0]    reg_psum_40_21;
wire signed[31:0]    reg_weight_40_22;
wire signed[31:0]    reg_psum_40_22;
wire signed[31:0]    reg_weight_40_23;
wire signed[31:0]    reg_psum_40_23;
wire signed[31:0]    reg_weight_40_24;
wire signed[31:0]    reg_psum_40_24;
wire signed[31:0]    reg_weight_40_25;
wire signed[31:0]    reg_psum_40_25;
wire signed[31:0]    reg_weight_40_26;
wire signed[31:0]    reg_psum_40_26;
wire signed[31:0]    reg_weight_40_27;
wire signed[31:0]    reg_psum_40_27;
wire signed[31:0]    reg_weight_40_28;
wire signed[31:0]    reg_psum_40_28;
wire signed[31:0]    reg_weight_40_29;
wire signed[31:0]    reg_psum_40_29;
wire signed[31:0]    reg_weight_40_30;
wire signed[31:0]    reg_psum_40_30;
wire signed[31:0]    reg_weight_40_31;
wire signed[31:0]    reg_psum_40_31;
wire signed[31:0]    reg_weight_40_32;
wire signed[31:0]    reg_psum_40_32;
wire signed[31:0]    reg_weight_40_33;
wire signed[31:0]    reg_psum_40_33;
wire signed[31:0]    reg_weight_40_34;
wire signed[31:0]    reg_psum_40_34;
wire signed[31:0]    reg_weight_40_35;
wire signed[31:0]    reg_psum_40_35;
wire signed[31:0]    reg_weight_40_36;
wire signed[31:0]    reg_psum_40_36;
wire signed[31:0]    reg_weight_40_37;
wire signed[31:0]    reg_psum_40_37;
wire signed[31:0]    reg_weight_40_38;
wire signed[31:0]    reg_psum_40_38;
wire signed[31:0]    reg_weight_40_39;
wire signed[31:0]    reg_psum_40_39;
wire signed[31:0]    reg_weight_40_40;
wire signed[31:0]    reg_psum_40_40;
wire signed[31:0]    reg_weight_40_41;
wire signed[31:0]    reg_psum_40_41;
wire signed[31:0]    reg_weight_40_42;
wire signed[31:0]    reg_psum_40_42;
wire signed[31:0]    reg_weight_40_43;
wire signed[31:0]    reg_psum_40_43;
wire signed[31:0]    reg_weight_40_44;
wire signed[31:0]    reg_psum_40_44;
wire signed[31:0]    reg_weight_40_45;
wire signed[31:0]    reg_psum_40_45;
wire signed[31:0]    reg_weight_40_46;
wire signed[31:0]    reg_psum_40_46;
wire signed[31:0]    reg_weight_40_47;
wire signed[31:0]    reg_psum_40_47;
wire signed[31:0]    reg_weight_40_48;
wire signed[31:0]    reg_psum_40_48;
wire signed[31:0]    reg_weight_40_49;
wire signed[31:0]    reg_psum_40_49;
wire signed[31:0]    reg_weight_40_50;
wire signed[31:0]    reg_psum_40_50;
wire signed[31:0]    reg_weight_40_51;
wire signed[31:0]    reg_psum_40_51;
wire signed[31:0]    reg_weight_40_52;
wire signed[31:0]    reg_psum_40_52;
wire signed[31:0]    reg_weight_40_53;
wire signed[31:0]    reg_psum_40_53;
wire signed[31:0]    reg_weight_40_54;
wire signed[31:0]    reg_psum_40_54;
wire signed[31:0]    reg_weight_40_55;
wire signed[31:0]    reg_psum_40_55;
wire signed[31:0]    reg_weight_40_56;
wire signed[31:0]    reg_psum_40_56;
wire signed[31:0]    reg_weight_40_57;
wire signed[31:0]    reg_psum_40_57;
wire signed[31:0]    reg_weight_40_58;
wire signed[31:0]    reg_psum_40_58;
wire signed[31:0]    reg_weight_40_59;
wire signed[31:0]    reg_psum_40_59;
wire signed[31:0]    reg_weight_40_60;
wire signed[31:0]    reg_psum_40_60;
wire signed[31:0]    reg_weight_40_61;
wire signed[31:0]    reg_psum_40_61;
wire signed[31:0]    reg_weight_40_62;
wire signed[31:0]    reg_psum_40_62;
wire signed[31:0]    reg_weight_40_63;
wire signed[31:0]    reg_psum_40_63;
wire signed[31:0]    reg_weight_41_0;
wire signed[31:0]    reg_psum_41_0;
wire signed[31:0]    reg_weight_41_1;
wire signed[31:0]    reg_psum_41_1;
wire signed[31:0]    reg_weight_41_2;
wire signed[31:0]    reg_psum_41_2;
wire signed[31:0]    reg_weight_41_3;
wire signed[31:0]    reg_psum_41_3;
wire signed[31:0]    reg_weight_41_4;
wire signed[31:0]    reg_psum_41_4;
wire signed[31:0]    reg_weight_41_5;
wire signed[31:0]    reg_psum_41_5;
wire signed[31:0]    reg_weight_41_6;
wire signed[31:0]    reg_psum_41_6;
wire signed[31:0]    reg_weight_41_7;
wire signed[31:0]    reg_psum_41_7;
wire signed[31:0]    reg_weight_41_8;
wire signed[31:0]    reg_psum_41_8;
wire signed[31:0]    reg_weight_41_9;
wire signed[31:0]    reg_psum_41_9;
wire signed[31:0]    reg_weight_41_10;
wire signed[31:0]    reg_psum_41_10;
wire signed[31:0]    reg_weight_41_11;
wire signed[31:0]    reg_psum_41_11;
wire signed[31:0]    reg_weight_41_12;
wire signed[31:0]    reg_psum_41_12;
wire signed[31:0]    reg_weight_41_13;
wire signed[31:0]    reg_psum_41_13;
wire signed[31:0]    reg_weight_41_14;
wire signed[31:0]    reg_psum_41_14;
wire signed[31:0]    reg_weight_41_15;
wire signed[31:0]    reg_psum_41_15;
wire signed[31:0]    reg_weight_41_16;
wire signed[31:0]    reg_psum_41_16;
wire signed[31:0]    reg_weight_41_17;
wire signed[31:0]    reg_psum_41_17;
wire signed[31:0]    reg_weight_41_18;
wire signed[31:0]    reg_psum_41_18;
wire signed[31:0]    reg_weight_41_19;
wire signed[31:0]    reg_psum_41_19;
wire signed[31:0]    reg_weight_41_20;
wire signed[31:0]    reg_psum_41_20;
wire signed[31:0]    reg_weight_41_21;
wire signed[31:0]    reg_psum_41_21;
wire signed[31:0]    reg_weight_41_22;
wire signed[31:0]    reg_psum_41_22;
wire signed[31:0]    reg_weight_41_23;
wire signed[31:0]    reg_psum_41_23;
wire signed[31:0]    reg_weight_41_24;
wire signed[31:0]    reg_psum_41_24;
wire signed[31:0]    reg_weight_41_25;
wire signed[31:0]    reg_psum_41_25;
wire signed[31:0]    reg_weight_41_26;
wire signed[31:0]    reg_psum_41_26;
wire signed[31:0]    reg_weight_41_27;
wire signed[31:0]    reg_psum_41_27;
wire signed[31:0]    reg_weight_41_28;
wire signed[31:0]    reg_psum_41_28;
wire signed[31:0]    reg_weight_41_29;
wire signed[31:0]    reg_psum_41_29;
wire signed[31:0]    reg_weight_41_30;
wire signed[31:0]    reg_psum_41_30;
wire signed[31:0]    reg_weight_41_31;
wire signed[31:0]    reg_psum_41_31;
wire signed[31:0]    reg_weight_41_32;
wire signed[31:0]    reg_psum_41_32;
wire signed[31:0]    reg_weight_41_33;
wire signed[31:0]    reg_psum_41_33;
wire signed[31:0]    reg_weight_41_34;
wire signed[31:0]    reg_psum_41_34;
wire signed[31:0]    reg_weight_41_35;
wire signed[31:0]    reg_psum_41_35;
wire signed[31:0]    reg_weight_41_36;
wire signed[31:0]    reg_psum_41_36;
wire signed[31:0]    reg_weight_41_37;
wire signed[31:0]    reg_psum_41_37;
wire signed[31:0]    reg_weight_41_38;
wire signed[31:0]    reg_psum_41_38;
wire signed[31:0]    reg_weight_41_39;
wire signed[31:0]    reg_psum_41_39;
wire signed[31:0]    reg_weight_41_40;
wire signed[31:0]    reg_psum_41_40;
wire signed[31:0]    reg_weight_41_41;
wire signed[31:0]    reg_psum_41_41;
wire signed[31:0]    reg_weight_41_42;
wire signed[31:0]    reg_psum_41_42;
wire signed[31:0]    reg_weight_41_43;
wire signed[31:0]    reg_psum_41_43;
wire signed[31:0]    reg_weight_41_44;
wire signed[31:0]    reg_psum_41_44;
wire signed[31:0]    reg_weight_41_45;
wire signed[31:0]    reg_psum_41_45;
wire signed[31:0]    reg_weight_41_46;
wire signed[31:0]    reg_psum_41_46;
wire signed[31:0]    reg_weight_41_47;
wire signed[31:0]    reg_psum_41_47;
wire signed[31:0]    reg_weight_41_48;
wire signed[31:0]    reg_psum_41_48;
wire signed[31:0]    reg_weight_41_49;
wire signed[31:0]    reg_psum_41_49;
wire signed[31:0]    reg_weight_41_50;
wire signed[31:0]    reg_psum_41_50;
wire signed[31:0]    reg_weight_41_51;
wire signed[31:0]    reg_psum_41_51;
wire signed[31:0]    reg_weight_41_52;
wire signed[31:0]    reg_psum_41_52;
wire signed[31:0]    reg_weight_41_53;
wire signed[31:0]    reg_psum_41_53;
wire signed[31:0]    reg_weight_41_54;
wire signed[31:0]    reg_psum_41_54;
wire signed[31:0]    reg_weight_41_55;
wire signed[31:0]    reg_psum_41_55;
wire signed[31:0]    reg_weight_41_56;
wire signed[31:0]    reg_psum_41_56;
wire signed[31:0]    reg_weight_41_57;
wire signed[31:0]    reg_psum_41_57;
wire signed[31:0]    reg_weight_41_58;
wire signed[31:0]    reg_psum_41_58;
wire signed[31:0]    reg_weight_41_59;
wire signed[31:0]    reg_psum_41_59;
wire signed[31:0]    reg_weight_41_60;
wire signed[31:0]    reg_psum_41_60;
wire signed[31:0]    reg_weight_41_61;
wire signed[31:0]    reg_psum_41_61;
wire signed[31:0]    reg_weight_41_62;
wire signed[31:0]    reg_psum_41_62;
wire signed[31:0]    reg_weight_41_63;
wire signed[31:0]    reg_psum_41_63;
wire signed[31:0]    reg_weight_42_0;
wire signed[31:0]    reg_psum_42_0;
wire signed[31:0]    reg_weight_42_1;
wire signed[31:0]    reg_psum_42_1;
wire signed[31:0]    reg_weight_42_2;
wire signed[31:0]    reg_psum_42_2;
wire signed[31:0]    reg_weight_42_3;
wire signed[31:0]    reg_psum_42_3;
wire signed[31:0]    reg_weight_42_4;
wire signed[31:0]    reg_psum_42_4;
wire signed[31:0]    reg_weight_42_5;
wire signed[31:0]    reg_psum_42_5;
wire signed[31:0]    reg_weight_42_6;
wire signed[31:0]    reg_psum_42_6;
wire signed[31:0]    reg_weight_42_7;
wire signed[31:0]    reg_psum_42_7;
wire signed[31:0]    reg_weight_42_8;
wire signed[31:0]    reg_psum_42_8;
wire signed[31:0]    reg_weight_42_9;
wire signed[31:0]    reg_psum_42_9;
wire signed[31:0]    reg_weight_42_10;
wire signed[31:0]    reg_psum_42_10;
wire signed[31:0]    reg_weight_42_11;
wire signed[31:0]    reg_psum_42_11;
wire signed[31:0]    reg_weight_42_12;
wire signed[31:0]    reg_psum_42_12;
wire signed[31:0]    reg_weight_42_13;
wire signed[31:0]    reg_psum_42_13;
wire signed[31:0]    reg_weight_42_14;
wire signed[31:0]    reg_psum_42_14;
wire signed[31:0]    reg_weight_42_15;
wire signed[31:0]    reg_psum_42_15;
wire signed[31:0]    reg_weight_42_16;
wire signed[31:0]    reg_psum_42_16;
wire signed[31:0]    reg_weight_42_17;
wire signed[31:0]    reg_psum_42_17;
wire signed[31:0]    reg_weight_42_18;
wire signed[31:0]    reg_psum_42_18;
wire signed[31:0]    reg_weight_42_19;
wire signed[31:0]    reg_psum_42_19;
wire signed[31:0]    reg_weight_42_20;
wire signed[31:0]    reg_psum_42_20;
wire signed[31:0]    reg_weight_42_21;
wire signed[31:0]    reg_psum_42_21;
wire signed[31:0]    reg_weight_42_22;
wire signed[31:0]    reg_psum_42_22;
wire signed[31:0]    reg_weight_42_23;
wire signed[31:0]    reg_psum_42_23;
wire signed[31:0]    reg_weight_42_24;
wire signed[31:0]    reg_psum_42_24;
wire signed[31:0]    reg_weight_42_25;
wire signed[31:0]    reg_psum_42_25;
wire signed[31:0]    reg_weight_42_26;
wire signed[31:0]    reg_psum_42_26;
wire signed[31:0]    reg_weight_42_27;
wire signed[31:0]    reg_psum_42_27;
wire signed[31:0]    reg_weight_42_28;
wire signed[31:0]    reg_psum_42_28;
wire signed[31:0]    reg_weight_42_29;
wire signed[31:0]    reg_psum_42_29;
wire signed[31:0]    reg_weight_42_30;
wire signed[31:0]    reg_psum_42_30;
wire signed[31:0]    reg_weight_42_31;
wire signed[31:0]    reg_psum_42_31;
wire signed[31:0]    reg_weight_42_32;
wire signed[31:0]    reg_psum_42_32;
wire signed[31:0]    reg_weight_42_33;
wire signed[31:0]    reg_psum_42_33;
wire signed[31:0]    reg_weight_42_34;
wire signed[31:0]    reg_psum_42_34;
wire signed[31:0]    reg_weight_42_35;
wire signed[31:0]    reg_psum_42_35;
wire signed[31:0]    reg_weight_42_36;
wire signed[31:0]    reg_psum_42_36;
wire signed[31:0]    reg_weight_42_37;
wire signed[31:0]    reg_psum_42_37;
wire signed[31:0]    reg_weight_42_38;
wire signed[31:0]    reg_psum_42_38;
wire signed[31:0]    reg_weight_42_39;
wire signed[31:0]    reg_psum_42_39;
wire signed[31:0]    reg_weight_42_40;
wire signed[31:0]    reg_psum_42_40;
wire signed[31:0]    reg_weight_42_41;
wire signed[31:0]    reg_psum_42_41;
wire signed[31:0]    reg_weight_42_42;
wire signed[31:0]    reg_psum_42_42;
wire signed[31:0]    reg_weight_42_43;
wire signed[31:0]    reg_psum_42_43;
wire signed[31:0]    reg_weight_42_44;
wire signed[31:0]    reg_psum_42_44;
wire signed[31:0]    reg_weight_42_45;
wire signed[31:0]    reg_psum_42_45;
wire signed[31:0]    reg_weight_42_46;
wire signed[31:0]    reg_psum_42_46;
wire signed[31:0]    reg_weight_42_47;
wire signed[31:0]    reg_psum_42_47;
wire signed[31:0]    reg_weight_42_48;
wire signed[31:0]    reg_psum_42_48;
wire signed[31:0]    reg_weight_42_49;
wire signed[31:0]    reg_psum_42_49;
wire signed[31:0]    reg_weight_42_50;
wire signed[31:0]    reg_psum_42_50;
wire signed[31:0]    reg_weight_42_51;
wire signed[31:0]    reg_psum_42_51;
wire signed[31:0]    reg_weight_42_52;
wire signed[31:0]    reg_psum_42_52;
wire signed[31:0]    reg_weight_42_53;
wire signed[31:0]    reg_psum_42_53;
wire signed[31:0]    reg_weight_42_54;
wire signed[31:0]    reg_psum_42_54;
wire signed[31:0]    reg_weight_42_55;
wire signed[31:0]    reg_psum_42_55;
wire signed[31:0]    reg_weight_42_56;
wire signed[31:0]    reg_psum_42_56;
wire signed[31:0]    reg_weight_42_57;
wire signed[31:0]    reg_psum_42_57;
wire signed[31:0]    reg_weight_42_58;
wire signed[31:0]    reg_psum_42_58;
wire signed[31:0]    reg_weight_42_59;
wire signed[31:0]    reg_psum_42_59;
wire signed[31:0]    reg_weight_42_60;
wire signed[31:0]    reg_psum_42_60;
wire signed[31:0]    reg_weight_42_61;
wire signed[31:0]    reg_psum_42_61;
wire signed[31:0]    reg_weight_42_62;
wire signed[31:0]    reg_psum_42_62;
wire signed[31:0]    reg_weight_42_63;
wire signed[31:0]    reg_psum_42_63;
wire signed[31:0]    reg_weight_43_0;
wire signed[31:0]    reg_psum_43_0;
wire signed[31:0]    reg_weight_43_1;
wire signed[31:0]    reg_psum_43_1;
wire signed[31:0]    reg_weight_43_2;
wire signed[31:0]    reg_psum_43_2;
wire signed[31:0]    reg_weight_43_3;
wire signed[31:0]    reg_psum_43_3;
wire signed[31:0]    reg_weight_43_4;
wire signed[31:0]    reg_psum_43_4;
wire signed[31:0]    reg_weight_43_5;
wire signed[31:0]    reg_psum_43_5;
wire signed[31:0]    reg_weight_43_6;
wire signed[31:0]    reg_psum_43_6;
wire signed[31:0]    reg_weight_43_7;
wire signed[31:0]    reg_psum_43_7;
wire signed[31:0]    reg_weight_43_8;
wire signed[31:0]    reg_psum_43_8;
wire signed[31:0]    reg_weight_43_9;
wire signed[31:0]    reg_psum_43_9;
wire signed[31:0]    reg_weight_43_10;
wire signed[31:0]    reg_psum_43_10;
wire signed[31:0]    reg_weight_43_11;
wire signed[31:0]    reg_psum_43_11;
wire signed[31:0]    reg_weight_43_12;
wire signed[31:0]    reg_psum_43_12;
wire signed[31:0]    reg_weight_43_13;
wire signed[31:0]    reg_psum_43_13;
wire signed[31:0]    reg_weight_43_14;
wire signed[31:0]    reg_psum_43_14;
wire signed[31:0]    reg_weight_43_15;
wire signed[31:0]    reg_psum_43_15;
wire signed[31:0]    reg_weight_43_16;
wire signed[31:0]    reg_psum_43_16;
wire signed[31:0]    reg_weight_43_17;
wire signed[31:0]    reg_psum_43_17;
wire signed[31:0]    reg_weight_43_18;
wire signed[31:0]    reg_psum_43_18;
wire signed[31:0]    reg_weight_43_19;
wire signed[31:0]    reg_psum_43_19;
wire signed[31:0]    reg_weight_43_20;
wire signed[31:0]    reg_psum_43_20;
wire signed[31:0]    reg_weight_43_21;
wire signed[31:0]    reg_psum_43_21;
wire signed[31:0]    reg_weight_43_22;
wire signed[31:0]    reg_psum_43_22;
wire signed[31:0]    reg_weight_43_23;
wire signed[31:0]    reg_psum_43_23;
wire signed[31:0]    reg_weight_43_24;
wire signed[31:0]    reg_psum_43_24;
wire signed[31:0]    reg_weight_43_25;
wire signed[31:0]    reg_psum_43_25;
wire signed[31:0]    reg_weight_43_26;
wire signed[31:0]    reg_psum_43_26;
wire signed[31:0]    reg_weight_43_27;
wire signed[31:0]    reg_psum_43_27;
wire signed[31:0]    reg_weight_43_28;
wire signed[31:0]    reg_psum_43_28;
wire signed[31:0]    reg_weight_43_29;
wire signed[31:0]    reg_psum_43_29;
wire signed[31:0]    reg_weight_43_30;
wire signed[31:0]    reg_psum_43_30;
wire signed[31:0]    reg_weight_43_31;
wire signed[31:0]    reg_psum_43_31;
wire signed[31:0]    reg_weight_43_32;
wire signed[31:0]    reg_psum_43_32;
wire signed[31:0]    reg_weight_43_33;
wire signed[31:0]    reg_psum_43_33;
wire signed[31:0]    reg_weight_43_34;
wire signed[31:0]    reg_psum_43_34;
wire signed[31:0]    reg_weight_43_35;
wire signed[31:0]    reg_psum_43_35;
wire signed[31:0]    reg_weight_43_36;
wire signed[31:0]    reg_psum_43_36;
wire signed[31:0]    reg_weight_43_37;
wire signed[31:0]    reg_psum_43_37;
wire signed[31:0]    reg_weight_43_38;
wire signed[31:0]    reg_psum_43_38;
wire signed[31:0]    reg_weight_43_39;
wire signed[31:0]    reg_psum_43_39;
wire signed[31:0]    reg_weight_43_40;
wire signed[31:0]    reg_psum_43_40;
wire signed[31:0]    reg_weight_43_41;
wire signed[31:0]    reg_psum_43_41;
wire signed[31:0]    reg_weight_43_42;
wire signed[31:0]    reg_psum_43_42;
wire signed[31:0]    reg_weight_43_43;
wire signed[31:0]    reg_psum_43_43;
wire signed[31:0]    reg_weight_43_44;
wire signed[31:0]    reg_psum_43_44;
wire signed[31:0]    reg_weight_43_45;
wire signed[31:0]    reg_psum_43_45;
wire signed[31:0]    reg_weight_43_46;
wire signed[31:0]    reg_psum_43_46;
wire signed[31:0]    reg_weight_43_47;
wire signed[31:0]    reg_psum_43_47;
wire signed[31:0]    reg_weight_43_48;
wire signed[31:0]    reg_psum_43_48;
wire signed[31:0]    reg_weight_43_49;
wire signed[31:0]    reg_psum_43_49;
wire signed[31:0]    reg_weight_43_50;
wire signed[31:0]    reg_psum_43_50;
wire signed[31:0]    reg_weight_43_51;
wire signed[31:0]    reg_psum_43_51;
wire signed[31:0]    reg_weight_43_52;
wire signed[31:0]    reg_psum_43_52;
wire signed[31:0]    reg_weight_43_53;
wire signed[31:0]    reg_psum_43_53;
wire signed[31:0]    reg_weight_43_54;
wire signed[31:0]    reg_psum_43_54;
wire signed[31:0]    reg_weight_43_55;
wire signed[31:0]    reg_psum_43_55;
wire signed[31:0]    reg_weight_43_56;
wire signed[31:0]    reg_psum_43_56;
wire signed[31:0]    reg_weight_43_57;
wire signed[31:0]    reg_psum_43_57;
wire signed[31:0]    reg_weight_43_58;
wire signed[31:0]    reg_psum_43_58;
wire signed[31:0]    reg_weight_43_59;
wire signed[31:0]    reg_psum_43_59;
wire signed[31:0]    reg_weight_43_60;
wire signed[31:0]    reg_psum_43_60;
wire signed[31:0]    reg_weight_43_61;
wire signed[31:0]    reg_psum_43_61;
wire signed[31:0]    reg_weight_43_62;
wire signed[31:0]    reg_psum_43_62;
wire signed[31:0]    reg_weight_43_63;
wire signed[31:0]    reg_psum_43_63;
wire signed[31:0]    reg_weight_44_0;
wire signed[31:0]    reg_psum_44_0;
wire signed[31:0]    reg_weight_44_1;
wire signed[31:0]    reg_psum_44_1;
wire signed[31:0]    reg_weight_44_2;
wire signed[31:0]    reg_psum_44_2;
wire signed[31:0]    reg_weight_44_3;
wire signed[31:0]    reg_psum_44_3;
wire signed[31:0]    reg_weight_44_4;
wire signed[31:0]    reg_psum_44_4;
wire signed[31:0]    reg_weight_44_5;
wire signed[31:0]    reg_psum_44_5;
wire signed[31:0]    reg_weight_44_6;
wire signed[31:0]    reg_psum_44_6;
wire signed[31:0]    reg_weight_44_7;
wire signed[31:0]    reg_psum_44_7;
wire signed[31:0]    reg_weight_44_8;
wire signed[31:0]    reg_psum_44_8;
wire signed[31:0]    reg_weight_44_9;
wire signed[31:0]    reg_psum_44_9;
wire signed[31:0]    reg_weight_44_10;
wire signed[31:0]    reg_psum_44_10;
wire signed[31:0]    reg_weight_44_11;
wire signed[31:0]    reg_psum_44_11;
wire signed[31:0]    reg_weight_44_12;
wire signed[31:0]    reg_psum_44_12;
wire signed[31:0]    reg_weight_44_13;
wire signed[31:0]    reg_psum_44_13;
wire signed[31:0]    reg_weight_44_14;
wire signed[31:0]    reg_psum_44_14;
wire signed[31:0]    reg_weight_44_15;
wire signed[31:0]    reg_psum_44_15;
wire signed[31:0]    reg_weight_44_16;
wire signed[31:0]    reg_psum_44_16;
wire signed[31:0]    reg_weight_44_17;
wire signed[31:0]    reg_psum_44_17;
wire signed[31:0]    reg_weight_44_18;
wire signed[31:0]    reg_psum_44_18;
wire signed[31:0]    reg_weight_44_19;
wire signed[31:0]    reg_psum_44_19;
wire signed[31:0]    reg_weight_44_20;
wire signed[31:0]    reg_psum_44_20;
wire signed[31:0]    reg_weight_44_21;
wire signed[31:0]    reg_psum_44_21;
wire signed[31:0]    reg_weight_44_22;
wire signed[31:0]    reg_psum_44_22;
wire signed[31:0]    reg_weight_44_23;
wire signed[31:0]    reg_psum_44_23;
wire signed[31:0]    reg_weight_44_24;
wire signed[31:0]    reg_psum_44_24;
wire signed[31:0]    reg_weight_44_25;
wire signed[31:0]    reg_psum_44_25;
wire signed[31:0]    reg_weight_44_26;
wire signed[31:0]    reg_psum_44_26;
wire signed[31:0]    reg_weight_44_27;
wire signed[31:0]    reg_psum_44_27;
wire signed[31:0]    reg_weight_44_28;
wire signed[31:0]    reg_psum_44_28;
wire signed[31:0]    reg_weight_44_29;
wire signed[31:0]    reg_psum_44_29;
wire signed[31:0]    reg_weight_44_30;
wire signed[31:0]    reg_psum_44_30;
wire signed[31:0]    reg_weight_44_31;
wire signed[31:0]    reg_psum_44_31;
wire signed[31:0]    reg_weight_44_32;
wire signed[31:0]    reg_psum_44_32;
wire signed[31:0]    reg_weight_44_33;
wire signed[31:0]    reg_psum_44_33;
wire signed[31:0]    reg_weight_44_34;
wire signed[31:0]    reg_psum_44_34;
wire signed[31:0]    reg_weight_44_35;
wire signed[31:0]    reg_psum_44_35;
wire signed[31:0]    reg_weight_44_36;
wire signed[31:0]    reg_psum_44_36;
wire signed[31:0]    reg_weight_44_37;
wire signed[31:0]    reg_psum_44_37;
wire signed[31:0]    reg_weight_44_38;
wire signed[31:0]    reg_psum_44_38;
wire signed[31:0]    reg_weight_44_39;
wire signed[31:0]    reg_psum_44_39;
wire signed[31:0]    reg_weight_44_40;
wire signed[31:0]    reg_psum_44_40;
wire signed[31:0]    reg_weight_44_41;
wire signed[31:0]    reg_psum_44_41;
wire signed[31:0]    reg_weight_44_42;
wire signed[31:0]    reg_psum_44_42;
wire signed[31:0]    reg_weight_44_43;
wire signed[31:0]    reg_psum_44_43;
wire signed[31:0]    reg_weight_44_44;
wire signed[31:0]    reg_psum_44_44;
wire signed[31:0]    reg_weight_44_45;
wire signed[31:0]    reg_psum_44_45;
wire signed[31:0]    reg_weight_44_46;
wire signed[31:0]    reg_psum_44_46;
wire signed[31:0]    reg_weight_44_47;
wire signed[31:0]    reg_psum_44_47;
wire signed[31:0]    reg_weight_44_48;
wire signed[31:0]    reg_psum_44_48;
wire signed[31:0]    reg_weight_44_49;
wire signed[31:0]    reg_psum_44_49;
wire signed[31:0]    reg_weight_44_50;
wire signed[31:0]    reg_psum_44_50;
wire signed[31:0]    reg_weight_44_51;
wire signed[31:0]    reg_psum_44_51;
wire signed[31:0]    reg_weight_44_52;
wire signed[31:0]    reg_psum_44_52;
wire signed[31:0]    reg_weight_44_53;
wire signed[31:0]    reg_psum_44_53;
wire signed[31:0]    reg_weight_44_54;
wire signed[31:0]    reg_psum_44_54;
wire signed[31:0]    reg_weight_44_55;
wire signed[31:0]    reg_psum_44_55;
wire signed[31:0]    reg_weight_44_56;
wire signed[31:0]    reg_psum_44_56;
wire signed[31:0]    reg_weight_44_57;
wire signed[31:0]    reg_psum_44_57;
wire signed[31:0]    reg_weight_44_58;
wire signed[31:0]    reg_psum_44_58;
wire signed[31:0]    reg_weight_44_59;
wire signed[31:0]    reg_psum_44_59;
wire signed[31:0]    reg_weight_44_60;
wire signed[31:0]    reg_psum_44_60;
wire signed[31:0]    reg_weight_44_61;
wire signed[31:0]    reg_psum_44_61;
wire signed[31:0]    reg_weight_44_62;
wire signed[31:0]    reg_psum_44_62;
wire signed[31:0]    reg_weight_44_63;
wire signed[31:0]    reg_psum_44_63;
wire signed[31:0]    reg_weight_45_0;
wire signed[31:0]    reg_psum_45_0;
wire signed[31:0]    reg_weight_45_1;
wire signed[31:0]    reg_psum_45_1;
wire signed[31:0]    reg_weight_45_2;
wire signed[31:0]    reg_psum_45_2;
wire signed[31:0]    reg_weight_45_3;
wire signed[31:0]    reg_psum_45_3;
wire signed[31:0]    reg_weight_45_4;
wire signed[31:0]    reg_psum_45_4;
wire signed[31:0]    reg_weight_45_5;
wire signed[31:0]    reg_psum_45_5;
wire signed[31:0]    reg_weight_45_6;
wire signed[31:0]    reg_psum_45_6;
wire signed[31:0]    reg_weight_45_7;
wire signed[31:0]    reg_psum_45_7;
wire signed[31:0]    reg_weight_45_8;
wire signed[31:0]    reg_psum_45_8;
wire signed[31:0]    reg_weight_45_9;
wire signed[31:0]    reg_psum_45_9;
wire signed[31:0]    reg_weight_45_10;
wire signed[31:0]    reg_psum_45_10;
wire signed[31:0]    reg_weight_45_11;
wire signed[31:0]    reg_psum_45_11;
wire signed[31:0]    reg_weight_45_12;
wire signed[31:0]    reg_psum_45_12;
wire signed[31:0]    reg_weight_45_13;
wire signed[31:0]    reg_psum_45_13;
wire signed[31:0]    reg_weight_45_14;
wire signed[31:0]    reg_psum_45_14;
wire signed[31:0]    reg_weight_45_15;
wire signed[31:0]    reg_psum_45_15;
wire signed[31:0]    reg_weight_45_16;
wire signed[31:0]    reg_psum_45_16;
wire signed[31:0]    reg_weight_45_17;
wire signed[31:0]    reg_psum_45_17;
wire signed[31:0]    reg_weight_45_18;
wire signed[31:0]    reg_psum_45_18;
wire signed[31:0]    reg_weight_45_19;
wire signed[31:0]    reg_psum_45_19;
wire signed[31:0]    reg_weight_45_20;
wire signed[31:0]    reg_psum_45_20;
wire signed[31:0]    reg_weight_45_21;
wire signed[31:0]    reg_psum_45_21;
wire signed[31:0]    reg_weight_45_22;
wire signed[31:0]    reg_psum_45_22;
wire signed[31:0]    reg_weight_45_23;
wire signed[31:0]    reg_psum_45_23;
wire signed[31:0]    reg_weight_45_24;
wire signed[31:0]    reg_psum_45_24;
wire signed[31:0]    reg_weight_45_25;
wire signed[31:0]    reg_psum_45_25;
wire signed[31:0]    reg_weight_45_26;
wire signed[31:0]    reg_psum_45_26;
wire signed[31:0]    reg_weight_45_27;
wire signed[31:0]    reg_psum_45_27;
wire signed[31:0]    reg_weight_45_28;
wire signed[31:0]    reg_psum_45_28;
wire signed[31:0]    reg_weight_45_29;
wire signed[31:0]    reg_psum_45_29;
wire signed[31:0]    reg_weight_45_30;
wire signed[31:0]    reg_psum_45_30;
wire signed[31:0]    reg_weight_45_31;
wire signed[31:0]    reg_psum_45_31;
wire signed[31:0]    reg_weight_45_32;
wire signed[31:0]    reg_psum_45_32;
wire signed[31:0]    reg_weight_45_33;
wire signed[31:0]    reg_psum_45_33;
wire signed[31:0]    reg_weight_45_34;
wire signed[31:0]    reg_psum_45_34;
wire signed[31:0]    reg_weight_45_35;
wire signed[31:0]    reg_psum_45_35;
wire signed[31:0]    reg_weight_45_36;
wire signed[31:0]    reg_psum_45_36;
wire signed[31:0]    reg_weight_45_37;
wire signed[31:0]    reg_psum_45_37;
wire signed[31:0]    reg_weight_45_38;
wire signed[31:0]    reg_psum_45_38;
wire signed[31:0]    reg_weight_45_39;
wire signed[31:0]    reg_psum_45_39;
wire signed[31:0]    reg_weight_45_40;
wire signed[31:0]    reg_psum_45_40;
wire signed[31:0]    reg_weight_45_41;
wire signed[31:0]    reg_psum_45_41;
wire signed[31:0]    reg_weight_45_42;
wire signed[31:0]    reg_psum_45_42;
wire signed[31:0]    reg_weight_45_43;
wire signed[31:0]    reg_psum_45_43;
wire signed[31:0]    reg_weight_45_44;
wire signed[31:0]    reg_psum_45_44;
wire signed[31:0]    reg_weight_45_45;
wire signed[31:0]    reg_psum_45_45;
wire signed[31:0]    reg_weight_45_46;
wire signed[31:0]    reg_psum_45_46;
wire signed[31:0]    reg_weight_45_47;
wire signed[31:0]    reg_psum_45_47;
wire signed[31:0]    reg_weight_45_48;
wire signed[31:0]    reg_psum_45_48;
wire signed[31:0]    reg_weight_45_49;
wire signed[31:0]    reg_psum_45_49;
wire signed[31:0]    reg_weight_45_50;
wire signed[31:0]    reg_psum_45_50;
wire signed[31:0]    reg_weight_45_51;
wire signed[31:0]    reg_psum_45_51;
wire signed[31:0]    reg_weight_45_52;
wire signed[31:0]    reg_psum_45_52;
wire signed[31:0]    reg_weight_45_53;
wire signed[31:0]    reg_psum_45_53;
wire signed[31:0]    reg_weight_45_54;
wire signed[31:0]    reg_psum_45_54;
wire signed[31:0]    reg_weight_45_55;
wire signed[31:0]    reg_psum_45_55;
wire signed[31:0]    reg_weight_45_56;
wire signed[31:0]    reg_psum_45_56;
wire signed[31:0]    reg_weight_45_57;
wire signed[31:0]    reg_psum_45_57;
wire signed[31:0]    reg_weight_45_58;
wire signed[31:0]    reg_psum_45_58;
wire signed[31:0]    reg_weight_45_59;
wire signed[31:0]    reg_psum_45_59;
wire signed[31:0]    reg_weight_45_60;
wire signed[31:0]    reg_psum_45_60;
wire signed[31:0]    reg_weight_45_61;
wire signed[31:0]    reg_psum_45_61;
wire signed[31:0]    reg_weight_45_62;
wire signed[31:0]    reg_psum_45_62;
wire signed[31:0]    reg_weight_45_63;
wire signed[31:0]    reg_psum_45_63;
wire signed[31:0]    reg_weight_46_0;
wire signed[31:0]    reg_psum_46_0;
wire signed[31:0]    reg_weight_46_1;
wire signed[31:0]    reg_psum_46_1;
wire signed[31:0]    reg_weight_46_2;
wire signed[31:0]    reg_psum_46_2;
wire signed[31:0]    reg_weight_46_3;
wire signed[31:0]    reg_psum_46_3;
wire signed[31:0]    reg_weight_46_4;
wire signed[31:0]    reg_psum_46_4;
wire signed[31:0]    reg_weight_46_5;
wire signed[31:0]    reg_psum_46_5;
wire signed[31:0]    reg_weight_46_6;
wire signed[31:0]    reg_psum_46_6;
wire signed[31:0]    reg_weight_46_7;
wire signed[31:0]    reg_psum_46_7;
wire signed[31:0]    reg_weight_46_8;
wire signed[31:0]    reg_psum_46_8;
wire signed[31:0]    reg_weight_46_9;
wire signed[31:0]    reg_psum_46_9;
wire signed[31:0]    reg_weight_46_10;
wire signed[31:0]    reg_psum_46_10;
wire signed[31:0]    reg_weight_46_11;
wire signed[31:0]    reg_psum_46_11;
wire signed[31:0]    reg_weight_46_12;
wire signed[31:0]    reg_psum_46_12;
wire signed[31:0]    reg_weight_46_13;
wire signed[31:0]    reg_psum_46_13;
wire signed[31:0]    reg_weight_46_14;
wire signed[31:0]    reg_psum_46_14;
wire signed[31:0]    reg_weight_46_15;
wire signed[31:0]    reg_psum_46_15;
wire signed[31:0]    reg_weight_46_16;
wire signed[31:0]    reg_psum_46_16;
wire signed[31:0]    reg_weight_46_17;
wire signed[31:0]    reg_psum_46_17;
wire signed[31:0]    reg_weight_46_18;
wire signed[31:0]    reg_psum_46_18;
wire signed[31:0]    reg_weight_46_19;
wire signed[31:0]    reg_psum_46_19;
wire signed[31:0]    reg_weight_46_20;
wire signed[31:0]    reg_psum_46_20;
wire signed[31:0]    reg_weight_46_21;
wire signed[31:0]    reg_psum_46_21;
wire signed[31:0]    reg_weight_46_22;
wire signed[31:0]    reg_psum_46_22;
wire signed[31:0]    reg_weight_46_23;
wire signed[31:0]    reg_psum_46_23;
wire signed[31:0]    reg_weight_46_24;
wire signed[31:0]    reg_psum_46_24;
wire signed[31:0]    reg_weight_46_25;
wire signed[31:0]    reg_psum_46_25;
wire signed[31:0]    reg_weight_46_26;
wire signed[31:0]    reg_psum_46_26;
wire signed[31:0]    reg_weight_46_27;
wire signed[31:0]    reg_psum_46_27;
wire signed[31:0]    reg_weight_46_28;
wire signed[31:0]    reg_psum_46_28;
wire signed[31:0]    reg_weight_46_29;
wire signed[31:0]    reg_psum_46_29;
wire signed[31:0]    reg_weight_46_30;
wire signed[31:0]    reg_psum_46_30;
wire signed[31:0]    reg_weight_46_31;
wire signed[31:0]    reg_psum_46_31;
wire signed[31:0]    reg_weight_46_32;
wire signed[31:0]    reg_psum_46_32;
wire signed[31:0]    reg_weight_46_33;
wire signed[31:0]    reg_psum_46_33;
wire signed[31:0]    reg_weight_46_34;
wire signed[31:0]    reg_psum_46_34;
wire signed[31:0]    reg_weight_46_35;
wire signed[31:0]    reg_psum_46_35;
wire signed[31:0]    reg_weight_46_36;
wire signed[31:0]    reg_psum_46_36;
wire signed[31:0]    reg_weight_46_37;
wire signed[31:0]    reg_psum_46_37;
wire signed[31:0]    reg_weight_46_38;
wire signed[31:0]    reg_psum_46_38;
wire signed[31:0]    reg_weight_46_39;
wire signed[31:0]    reg_psum_46_39;
wire signed[31:0]    reg_weight_46_40;
wire signed[31:0]    reg_psum_46_40;
wire signed[31:0]    reg_weight_46_41;
wire signed[31:0]    reg_psum_46_41;
wire signed[31:0]    reg_weight_46_42;
wire signed[31:0]    reg_psum_46_42;
wire signed[31:0]    reg_weight_46_43;
wire signed[31:0]    reg_psum_46_43;
wire signed[31:0]    reg_weight_46_44;
wire signed[31:0]    reg_psum_46_44;
wire signed[31:0]    reg_weight_46_45;
wire signed[31:0]    reg_psum_46_45;
wire signed[31:0]    reg_weight_46_46;
wire signed[31:0]    reg_psum_46_46;
wire signed[31:0]    reg_weight_46_47;
wire signed[31:0]    reg_psum_46_47;
wire signed[31:0]    reg_weight_46_48;
wire signed[31:0]    reg_psum_46_48;
wire signed[31:0]    reg_weight_46_49;
wire signed[31:0]    reg_psum_46_49;
wire signed[31:0]    reg_weight_46_50;
wire signed[31:0]    reg_psum_46_50;
wire signed[31:0]    reg_weight_46_51;
wire signed[31:0]    reg_psum_46_51;
wire signed[31:0]    reg_weight_46_52;
wire signed[31:0]    reg_psum_46_52;
wire signed[31:0]    reg_weight_46_53;
wire signed[31:0]    reg_psum_46_53;
wire signed[31:0]    reg_weight_46_54;
wire signed[31:0]    reg_psum_46_54;
wire signed[31:0]    reg_weight_46_55;
wire signed[31:0]    reg_psum_46_55;
wire signed[31:0]    reg_weight_46_56;
wire signed[31:0]    reg_psum_46_56;
wire signed[31:0]    reg_weight_46_57;
wire signed[31:0]    reg_psum_46_57;
wire signed[31:0]    reg_weight_46_58;
wire signed[31:0]    reg_psum_46_58;
wire signed[31:0]    reg_weight_46_59;
wire signed[31:0]    reg_psum_46_59;
wire signed[31:0]    reg_weight_46_60;
wire signed[31:0]    reg_psum_46_60;
wire signed[31:0]    reg_weight_46_61;
wire signed[31:0]    reg_psum_46_61;
wire signed[31:0]    reg_weight_46_62;
wire signed[31:0]    reg_psum_46_62;
wire signed[31:0]    reg_weight_46_63;
wire signed[31:0]    reg_psum_46_63;
wire signed[31:0]    reg_weight_47_0;
wire signed[31:0]    reg_psum_47_0;
wire signed[31:0]    reg_weight_47_1;
wire signed[31:0]    reg_psum_47_1;
wire signed[31:0]    reg_weight_47_2;
wire signed[31:0]    reg_psum_47_2;
wire signed[31:0]    reg_weight_47_3;
wire signed[31:0]    reg_psum_47_3;
wire signed[31:0]    reg_weight_47_4;
wire signed[31:0]    reg_psum_47_4;
wire signed[31:0]    reg_weight_47_5;
wire signed[31:0]    reg_psum_47_5;
wire signed[31:0]    reg_weight_47_6;
wire signed[31:0]    reg_psum_47_6;
wire signed[31:0]    reg_weight_47_7;
wire signed[31:0]    reg_psum_47_7;
wire signed[31:0]    reg_weight_47_8;
wire signed[31:0]    reg_psum_47_8;
wire signed[31:0]    reg_weight_47_9;
wire signed[31:0]    reg_psum_47_9;
wire signed[31:0]    reg_weight_47_10;
wire signed[31:0]    reg_psum_47_10;
wire signed[31:0]    reg_weight_47_11;
wire signed[31:0]    reg_psum_47_11;
wire signed[31:0]    reg_weight_47_12;
wire signed[31:0]    reg_psum_47_12;
wire signed[31:0]    reg_weight_47_13;
wire signed[31:0]    reg_psum_47_13;
wire signed[31:0]    reg_weight_47_14;
wire signed[31:0]    reg_psum_47_14;
wire signed[31:0]    reg_weight_47_15;
wire signed[31:0]    reg_psum_47_15;
wire signed[31:0]    reg_weight_47_16;
wire signed[31:0]    reg_psum_47_16;
wire signed[31:0]    reg_weight_47_17;
wire signed[31:0]    reg_psum_47_17;
wire signed[31:0]    reg_weight_47_18;
wire signed[31:0]    reg_psum_47_18;
wire signed[31:0]    reg_weight_47_19;
wire signed[31:0]    reg_psum_47_19;
wire signed[31:0]    reg_weight_47_20;
wire signed[31:0]    reg_psum_47_20;
wire signed[31:0]    reg_weight_47_21;
wire signed[31:0]    reg_psum_47_21;
wire signed[31:0]    reg_weight_47_22;
wire signed[31:0]    reg_psum_47_22;
wire signed[31:0]    reg_weight_47_23;
wire signed[31:0]    reg_psum_47_23;
wire signed[31:0]    reg_weight_47_24;
wire signed[31:0]    reg_psum_47_24;
wire signed[31:0]    reg_weight_47_25;
wire signed[31:0]    reg_psum_47_25;
wire signed[31:0]    reg_weight_47_26;
wire signed[31:0]    reg_psum_47_26;
wire signed[31:0]    reg_weight_47_27;
wire signed[31:0]    reg_psum_47_27;
wire signed[31:0]    reg_weight_47_28;
wire signed[31:0]    reg_psum_47_28;
wire signed[31:0]    reg_weight_47_29;
wire signed[31:0]    reg_psum_47_29;
wire signed[31:0]    reg_weight_47_30;
wire signed[31:0]    reg_psum_47_30;
wire signed[31:0]    reg_weight_47_31;
wire signed[31:0]    reg_psum_47_31;
wire signed[31:0]    reg_weight_47_32;
wire signed[31:0]    reg_psum_47_32;
wire signed[31:0]    reg_weight_47_33;
wire signed[31:0]    reg_psum_47_33;
wire signed[31:0]    reg_weight_47_34;
wire signed[31:0]    reg_psum_47_34;
wire signed[31:0]    reg_weight_47_35;
wire signed[31:0]    reg_psum_47_35;
wire signed[31:0]    reg_weight_47_36;
wire signed[31:0]    reg_psum_47_36;
wire signed[31:0]    reg_weight_47_37;
wire signed[31:0]    reg_psum_47_37;
wire signed[31:0]    reg_weight_47_38;
wire signed[31:0]    reg_psum_47_38;
wire signed[31:0]    reg_weight_47_39;
wire signed[31:0]    reg_psum_47_39;
wire signed[31:0]    reg_weight_47_40;
wire signed[31:0]    reg_psum_47_40;
wire signed[31:0]    reg_weight_47_41;
wire signed[31:0]    reg_psum_47_41;
wire signed[31:0]    reg_weight_47_42;
wire signed[31:0]    reg_psum_47_42;
wire signed[31:0]    reg_weight_47_43;
wire signed[31:0]    reg_psum_47_43;
wire signed[31:0]    reg_weight_47_44;
wire signed[31:0]    reg_psum_47_44;
wire signed[31:0]    reg_weight_47_45;
wire signed[31:0]    reg_psum_47_45;
wire signed[31:0]    reg_weight_47_46;
wire signed[31:0]    reg_psum_47_46;
wire signed[31:0]    reg_weight_47_47;
wire signed[31:0]    reg_psum_47_47;
wire signed[31:0]    reg_weight_47_48;
wire signed[31:0]    reg_psum_47_48;
wire signed[31:0]    reg_weight_47_49;
wire signed[31:0]    reg_psum_47_49;
wire signed[31:0]    reg_weight_47_50;
wire signed[31:0]    reg_psum_47_50;
wire signed[31:0]    reg_weight_47_51;
wire signed[31:0]    reg_psum_47_51;
wire signed[31:0]    reg_weight_47_52;
wire signed[31:0]    reg_psum_47_52;
wire signed[31:0]    reg_weight_47_53;
wire signed[31:0]    reg_psum_47_53;
wire signed[31:0]    reg_weight_47_54;
wire signed[31:0]    reg_psum_47_54;
wire signed[31:0]    reg_weight_47_55;
wire signed[31:0]    reg_psum_47_55;
wire signed[31:0]    reg_weight_47_56;
wire signed[31:0]    reg_psum_47_56;
wire signed[31:0]    reg_weight_47_57;
wire signed[31:0]    reg_psum_47_57;
wire signed[31:0]    reg_weight_47_58;
wire signed[31:0]    reg_psum_47_58;
wire signed[31:0]    reg_weight_47_59;
wire signed[31:0]    reg_psum_47_59;
wire signed[31:0]    reg_weight_47_60;
wire signed[31:0]    reg_psum_47_60;
wire signed[31:0]    reg_weight_47_61;
wire signed[31:0]    reg_psum_47_61;
wire signed[31:0]    reg_weight_47_62;
wire signed[31:0]    reg_psum_47_62;
wire signed[31:0]    reg_weight_47_63;
wire signed[31:0]    reg_psum_47_63;
wire signed[31:0]    reg_weight_48_0;
wire signed[31:0]    reg_psum_48_0;
wire signed[31:0]    reg_weight_48_1;
wire signed[31:0]    reg_psum_48_1;
wire signed[31:0]    reg_weight_48_2;
wire signed[31:0]    reg_psum_48_2;
wire signed[31:0]    reg_weight_48_3;
wire signed[31:0]    reg_psum_48_3;
wire signed[31:0]    reg_weight_48_4;
wire signed[31:0]    reg_psum_48_4;
wire signed[31:0]    reg_weight_48_5;
wire signed[31:0]    reg_psum_48_5;
wire signed[31:0]    reg_weight_48_6;
wire signed[31:0]    reg_psum_48_6;
wire signed[31:0]    reg_weight_48_7;
wire signed[31:0]    reg_psum_48_7;
wire signed[31:0]    reg_weight_48_8;
wire signed[31:0]    reg_psum_48_8;
wire signed[31:0]    reg_weight_48_9;
wire signed[31:0]    reg_psum_48_9;
wire signed[31:0]    reg_weight_48_10;
wire signed[31:0]    reg_psum_48_10;
wire signed[31:0]    reg_weight_48_11;
wire signed[31:0]    reg_psum_48_11;
wire signed[31:0]    reg_weight_48_12;
wire signed[31:0]    reg_psum_48_12;
wire signed[31:0]    reg_weight_48_13;
wire signed[31:0]    reg_psum_48_13;
wire signed[31:0]    reg_weight_48_14;
wire signed[31:0]    reg_psum_48_14;
wire signed[31:0]    reg_weight_48_15;
wire signed[31:0]    reg_psum_48_15;
wire signed[31:0]    reg_weight_48_16;
wire signed[31:0]    reg_psum_48_16;
wire signed[31:0]    reg_weight_48_17;
wire signed[31:0]    reg_psum_48_17;
wire signed[31:0]    reg_weight_48_18;
wire signed[31:0]    reg_psum_48_18;
wire signed[31:0]    reg_weight_48_19;
wire signed[31:0]    reg_psum_48_19;
wire signed[31:0]    reg_weight_48_20;
wire signed[31:0]    reg_psum_48_20;
wire signed[31:0]    reg_weight_48_21;
wire signed[31:0]    reg_psum_48_21;
wire signed[31:0]    reg_weight_48_22;
wire signed[31:0]    reg_psum_48_22;
wire signed[31:0]    reg_weight_48_23;
wire signed[31:0]    reg_psum_48_23;
wire signed[31:0]    reg_weight_48_24;
wire signed[31:0]    reg_psum_48_24;
wire signed[31:0]    reg_weight_48_25;
wire signed[31:0]    reg_psum_48_25;
wire signed[31:0]    reg_weight_48_26;
wire signed[31:0]    reg_psum_48_26;
wire signed[31:0]    reg_weight_48_27;
wire signed[31:0]    reg_psum_48_27;
wire signed[31:0]    reg_weight_48_28;
wire signed[31:0]    reg_psum_48_28;
wire signed[31:0]    reg_weight_48_29;
wire signed[31:0]    reg_psum_48_29;
wire signed[31:0]    reg_weight_48_30;
wire signed[31:0]    reg_psum_48_30;
wire signed[31:0]    reg_weight_48_31;
wire signed[31:0]    reg_psum_48_31;
wire signed[31:0]    reg_weight_48_32;
wire signed[31:0]    reg_psum_48_32;
wire signed[31:0]    reg_weight_48_33;
wire signed[31:0]    reg_psum_48_33;
wire signed[31:0]    reg_weight_48_34;
wire signed[31:0]    reg_psum_48_34;
wire signed[31:0]    reg_weight_48_35;
wire signed[31:0]    reg_psum_48_35;
wire signed[31:0]    reg_weight_48_36;
wire signed[31:0]    reg_psum_48_36;
wire signed[31:0]    reg_weight_48_37;
wire signed[31:0]    reg_psum_48_37;
wire signed[31:0]    reg_weight_48_38;
wire signed[31:0]    reg_psum_48_38;
wire signed[31:0]    reg_weight_48_39;
wire signed[31:0]    reg_psum_48_39;
wire signed[31:0]    reg_weight_48_40;
wire signed[31:0]    reg_psum_48_40;
wire signed[31:0]    reg_weight_48_41;
wire signed[31:0]    reg_psum_48_41;
wire signed[31:0]    reg_weight_48_42;
wire signed[31:0]    reg_psum_48_42;
wire signed[31:0]    reg_weight_48_43;
wire signed[31:0]    reg_psum_48_43;
wire signed[31:0]    reg_weight_48_44;
wire signed[31:0]    reg_psum_48_44;
wire signed[31:0]    reg_weight_48_45;
wire signed[31:0]    reg_psum_48_45;
wire signed[31:0]    reg_weight_48_46;
wire signed[31:0]    reg_psum_48_46;
wire signed[31:0]    reg_weight_48_47;
wire signed[31:0]    reg_psum_48_47;
wire signed[31:0]    reg_weight_48_48;
wire signed[31:0]    reg_psum_48_48;
wire signed[31:0]    reg_weight_48_49;
wire signed[31:0]    reg_psum_48_49;
wire signed[31:0]    reg_weight_48_50;
wire signed[31:0]    reg_psum_48_50;
wire signed[31:0]    reg_weight_48_51;
wire signed[31:0]    reg_psum_48_51;
wire signed[31:0]    reg_weight_48_52;
wire signed[31:0]    reg_psum_48_52;
wire signed[31:0]    reg_weight_48_53;
wire signed[31:0]    reg_psum_48_53;
wire signed[31:0]    reg_weight_48_54;
wire signed[31:0]    reg_psum_48_54;
wire signed[31:0]    reg_weight_48_55;
wire signed[31:0]    reg_psum_48_55;
wire signed[31:0]    reg_weight_48_56;
wire signed[31:0]    reg_psum_48_56;
wire signed[31:0]    reg_weight_48_57;
wire signed[31:0]    reg_psum_48_57;
wire signed[31:0]    reg_weight_48_58;
wire signed[31:0]    reg_psum_48_58;
wire signed[31:0]    reg_weight_48_59;
wire signed[31:0]    reg_psum_48_59;
wire signed[31:0]    reg_weight_48_60;
wire signed[31:0]    reg_psum_48_60;
wire signed[31:0]    reg_weight_48_61;
wire signed[31:0]    reg_psum_48_61;
wire signed[31:0]    reg_weight_48_62;
wire signed[31:0]    reg_psum_48_62;
wire signed[31:0]    reg_weight_48_63;
wire signed[31:0]    reg_psum_48_63;
wire signed[31:0]    reg_weight_49_0;
wire signed[31:0]    reg_psum_49_0;
wire signed[31:0]    reg_weight_49_1;
wire signed[31:0]    reg_psum_49_1;
wire signed[31:0]    reg_weight_49_2;
wire signed[31:0]    reg_psum_49_2;
wire signed[31:0]    reg_weight_49_3;
wire signed[31:0]    reg_psum_49_3;
wire signed[31:0]    reg_weight_49_4;
wire signed[31:0]    reg_psum_49_4;
wire signed[31:0]    reg_weight_49_5;
wire signed[31:0]    reg_psum_49_5;
wire signed[31:0]    reg_weight_49_6;
wire signed[31:0]    reg_psum_49_6;
wire signed[31:0]    reg_weight_49_7;
wire signed[31:0]    reg_psum_49_7;
wire signed[31:0]    reg_weight_49_8;
wire signed[31:0]    reg_psum_49_8;
wire signed[31:0]    reg_weight_49_9;
wire signed[31:0]    reg_psum_49_9;
wire signed[31:0]    reg_weight_49_10;
wire signed[31:0]    reg_psum_49_10;
wire signed[31:0]    reg_weight_49_11;
wire signed[31:0]    reg_psum_49_11;
wire signed[31:0]    reg_weight_49_12;
wire signed[31:0]    reg_psum_49_12;
wire signed[31:0]    reg_weight_49_13;
wire signed[31:0]    reg_psum_49_13;
wire signed[31:0]    reg_weight_49_14;
wire signed[31:0]    reg_psum_49_14;
wire signed[31:0]    reg_weight_49_15;
wire signed[31:0]    reg_psum_49_15;
wire signed[31:0]    reg_weight_49_16;
wire signed[31:0]    reg_psum_49_16;
wire signed[31:0]    reg_weight_49_17;
wire signed[31:0]    reg_psum_49_17;
wire signed[31:0]    reg_weight_49_18;
wire signed[31:0]    reg_psum_49_18;
wire signed[31:0]    reg_weight_49_19;
wire signed[31:0]    reg_psum_49_19;
wire signed[31:0]    reg_weight_49_20;
wire signed[31:0]    reg_psum_49_20;
wire signed[31:0]    reg_weight_49_21;
wire signed[31:0]    reg_psum_49_21;
wire signed[31:0]    reg_weight_49_22;
wire signed[31:0]    reg_psum_49_22;
wire signed[31:0]    reg_weight_49_23;
wire signed[31:0]    reg_psum_49_23;
wire signed[31:0]    reg_weight_49_24;
wire signed[31:0]    reg_psum_49_24;
wire signed[31:0]    reg_weight_49_25;
wire signed[31:0]    reg_psum_49_25;
wire signed[31:0]    reg_weight_49_26;
wire signed[31:0]    reg_psum_49_26;
wire signed[31:0]    reg_weight_49_27;
wire signed[31:0]    reg_psum_49_27;
wire signed[31:0]    reg_weight_49_28;
wire signed[31:0]    reg_psum_49_28;
wire signed[31:0]    reg_weight_49_29;
wire signed[31:0]    reg_psum_49_29;
wire signed[31:0]    reg_weight_49_30;
wire signed[31:0]    reg_psum_49_30;
wire signed[31:0]    reg_weight_49_31;
wire signed[31:0]    reg_psum_49_31;
wire signed[31:0]    reg_weight_49_32;
wire signed[31:0]    reg_psum_49_32;
wire signed[31:0]    reg_weight_49_33;
wire signed[31:0]    reg_psum_49_33;
wire signed[31:0]    reg_weight_49_34;
wire signed[31:0]    reg_psum_49_34;
wire signed[31:0]    reg_weight_49_35;
wire signed[31:0]    reg_psum_49_35;
wire signed[31:0]    reg_weight_49_36;
wire signed[31:0]    reg_psum_49_36;
wire signed[31:0]    reg_weight_49_37;
wire signed[31:0]    reg_psum_49_37;
wire signed[31:0]    reg_weight_49_38;
wire signed[31:0]    reg_psum_49_38;
wire signed[31:0]    reg_weight_49_39;
wire signed[31:0]    reg_psum_49_39;
wire signed[31:0]    reg_weight_49_40;
wire signed[31:0]    reg_psum_49_40;
wire signed[31:0]    reg_weight_49_41;
wire signed[31:0]    reg_psum_49_41;
wire signed[31:0]    reg_weight_49_42;
wire signed[31:0]    reg_psum_49_42;
wire signed[31:0]    reg_weight_49_43;
wire signed[31:0]    reg_psum_49_43;
wire signed[31:0]    reg_weight_49_44;
wire signed[31:0]    reg_psum_49_44;
wire signed[31:0]    reg_weight_49_45;
wire signed[31:0]    reg_psum_49_45;
wire signed[31:0]    reg_weight_49_46;
wire signed[31:0]    reg_psum_49_46;
wire signed[31:0]    reg_weight_49_47;
wire signed[31:0]    reg_psum_49_47;
wire signed[31:0]    reg_weight_49_48;
wire signed[31:0]    reg_psum_49_48;
wire signed[31:0]    reg_weight_49_49;
wire signed[31:0]    reg_psum_49_49;
wire signed[31:0]    reg_weight_49_50;
wire signed[31:0]    reg_psum_49_50;
wire signed[31:0]    reg_weight_49_51;
wire signed[31:0]    reg_psum_49_51;
wire signed[31:0]    reg_weight_49_52;
wire signed[31:0]    reg_psum_49_52;
wire signed[31:0]    reg_weight_49_53;
wire signed[31:0]    reg_psum_49_53;
wire signed[31:0]    reg_weight_49_54;
wire signed[31:0]    reg_psum_49_54;
wire signed[31:0]    reg_weight_49_55;
wire signed[31:0]    reg_psum_49_55;
wire signed[31:0]    reg_weight_49_56;
wire signed[31:0]    reg_psum_49_56;
wire signed[31:0]    reg_weight_49_57;
wire signed[31:0]    reg_psum_49_57;
wire signed[31:0]    reg_weight_49_58;
wire signed[31:0]    reg_psum_49_58;
wire signed[31:0]    reg_weight_49_59;
wire signed[31:0]    reg_psum_49_59;
wire signed[31:0]    reg_weight_49_60;
wire signed[31:0]    reg_psum_49_60;
wire signed[31:0]    reg_weight_49_61;
wire signed[31:0]    reg_psum_49_61;
wire signed[31:0]    reg_weight_49_62;
wire signed[31:0]    reg_psum_49_62;
wire signed[31:0]    reg_weight_49_63;
wire signed[31:0]    reg_psum_49_63;
wire signed[31:0]    reg_weight_50_0;
wire signed[31:0]    reg_psum_50_0;
wire signed[31:0]    reg_weight_50_1;
wire signed[31:0]    reg_psum_50_1;
wire signed[31:0]    reg_weight_50_2;
wire signed[31:0]    reg_psum_50_2;
wire signed[31:0]    reg_weight_50_3;
wire signed[31:0]    reg_psum_50_3;
wire signed[31:0]    reg_weight_50_4;
wire signed[31:0]    reg_psum_50_4;
wire signed[31:0]    reg_weight_50_5;
wire signed[31:0]    reg_psum_50_5;
wire signed[31:0]    reg_weight_50_6;
wire signed[31:0]    reg_psum_50_6;
wire signed[31:0]    reg_weight_50_7;
wire signed[31:0]    reg_psum_50_7;
wire signed[31:0]    reg_weight_50_8;
wire signed[31:0]    reg_psum_50_8;
wire signed[31:0]    reg_weight_50_9;
wire signed[31:0]    reg_psum_50_9;
wire signed[31:0]    reg_weight_50_10;
wire signed[31:0]    reg_psum_50_10;
wire signed[31:0]    reg_weight_50_11;
wire signed[31:0]    reg_psum_50_11;
wire signed[31:0]    reg_weight_50_12;
wire signed[31:0]    reg_psum_50_12;
wire signed[31:0]    reg_weight_50_13;
wire signed[31:0]    reg_psum_50_13;
wire signed[31:0]    reg_weight_50_14;
wire signed[31:0]    reg_psum_50_14;
wire signed[31:0]    reg_weight_50_15;
wire signed[31:0]    reg_psum_50_15;
wire signed[31:0]    reg_weight_50_16;
wire signed[31:0]    reg_psum_50_16;
wire signed[31:0]    reg_weight_50_17;
wire signed[31:0]    reg_psum_50_17;
wire signed[31:0]    reg_weight_50_18;
wire signed[31:0]    reg_psum_50_18;
wire signed[31:0]    reg_weight_50_19;
wire signed[31:0]    reg_psum_50_19;
wire signed[31:0]    reg_weight_50_20;
wire signed[31:0]    reg_psum_50_20;
wire signed[31:0]    reg_weight_50_21;
wire signed[31:0]    reg_psum_50_21;
wire signed[31:0]    reg_weight_50_22;
wire signed[31:0]    reg_psum_50_22;
wire signed[31:0]    reg_weight_50_23;
wire signed[31:0]    reg_psum_50_23;
wire signed[31:0]    reg_weight_50_24;
wire signed[31:0]    reg_psum_50_24;
wire signed[31:0]    reg_weight_50_25;
wire signed[31:0]    reg_psum_50_25;
wire signed[31:0]    reg_weight_50_26;
wire signed[31:0]    reg_psum_50_26;
wire signed[31:0]    reg_weight_50_27;
wire signed[31:0]    reg_psum_50_27;
wire signed[31:0]    reg_weight_50_28;
wire signed[31:0]    reg_psum_50_28;
wire signed[31:0]    reg_weight_50_29;
wire signed[31:0]    reg_psum_50_29;
wire signed[31:0]    reg_weight_50_30;
wire signed[31:0]    reg_psum_50_30;
wire signed[31:0]    reg_weight_50_31;
wire signed[31:0]    reg_psum_50_31;
wire signed[31:0]    reg_weight_50_32;
wire signed[31:0]    reg_psum_50_32;
wire signed[31:0]    reg_weight_50_33;
wire signed[31:0]    reg_psum_50_33;
wire signed[31:0]    reg_weight_50_34;
wire signed[31:0]    reg_psum_50_34;
wire signed[31:0]    reg_weight_50_35;
wire signed[31:0]    reg_psum_50_35;
wire signed[31:0]    reg_weight_50_36;
wire signed[31:0]    reg_psum_50_36;
wire signed[31:0]    reg_weight_50_37;
wire signed[31:0]    reg_psum_50_37;
wire signed[31:0]    reg_weight_50_38;
wire signed[31:0]    reg_psum_50_38;
wire signed[31:0]    reg_weight_50_39;
wire signed[31:0]    reg_psum_50_39;
wire signed[31:0]    reg_weight_50_40;
wire signed[31:0]    reg_psum_50_40;
wire signed[31:0]    reg_weight_50_41;
wire signed[31:0]    reg_psum_50_41;
wire signed[31:0]    reg_weight_50_42;
wire signed[31:0]    reg_psum_50_42;
wire signed[31:0]    reg_weight_50_43;
wire signed[31:0]    reg_psum_50_43;
wire signed[31:0]    reg_weight_50_44;
wire signed[31:0]    reg_psum_50_44;
wire signed[31:0]    reg_weight_50_45;
wire signed[31:0]    reg_psum_50_45;
wire signed[31:0]    reg_weight_50_46;
wire signed[31:0]    reg_psum_50_46;
wire signed[31:0]    reg_weight_50_47;
wire signed[31:0]    reg_psum_50_47;
wire signed[31:0]    reg_weight_50_48;
wire signed[31:0]    reg_psum_50_48;
wire signed[31:0]    reg_weight_50_49;
wire signed[31:0]    reg_psum_50_49;
wire signed[31:0]    reg_weight_50_50;
wire signed[31:0]    reg_psum_50_50;
wire signed[31:0]    reg_weight_50_51;
wire signed[31:0]    reg_psum_50_51;
wire signed[31:0]    reg_weight_50_52;
wire signed[31:0]    reg_psum_50_52;
wire signed[31:0]    reg_weight_50_53;
wire signed[31:0]    reg_psum_50_53;
wire signed[31:0]    reg_weight_50_54;
wire signed[31:0]    reg_psum_50_54;
wire signed[31:0]    reg_weight_50_55;
wire signed[31:0]    reg_psum_50_55;
wire signed[31:0]    reg_weight_50_56;
wire signed[31:0]    reg_psum_50_56;
wire signed[31:0]    reg_weight_50_57;
wire signed[31:0]    reg_psum_50_57;
wire signed[31:0]    reg_weight_50_58;
wire signed[31:0]    reg_psum_50_58;
wire signed[31:0]    reg_weight_50_59;
wire signed[31:0]    reg_psum_50_59;
wire signed[31:0]    reg_weight_50_60;
wire signed[31:0]    reg_psum_50_60;
wire signed[31:0]    reg_weight_50_61;
wire signed[31:0]    reg_psum_50_61;
wire signed[31:0]    reg_weight_50_62;
wire signed[31:0]    reg_psum_50_62;
wire signed[31:0]    reg_weight_50_63;
wire signed[31:0]    reg_psum_50_63;
wire signed[31:0]    reg_weight_51_0;
wire signed[31:0]    reg_psum_51_0;
wire signed[31:0]    reg_weight_51_1;
wire signed[31:0]    reg_psum_51_1;
wire signed[31:0]    reg_weight_51_2;
wire signed[31:0]    reg_psum_51_2;
wire signed[31:0]    reg_weight_51_3;
wire signed[31:0]    reg_psum_51_3;
wire signed[31:0]    reg_weight_51_4;
wire signed[31:0]    reg_psum_51_4;
wire signed[31:0]    reg_weight_51_5;
wire signed[31:0]    reg_psum_51_5;
wire signed[31:0]    reg_weight_51_6;
wire signed[31:0]    reg_psum_51_6;
wire signed[31:0]    reg_weight_51_7;
wire signed[31:0]    reg_psum_51_7;
wire signed[31:0]    reg_weight_51_8;
wire signed[31:0]    reg_psum_51_8;
wire signed[31:0]    reg_weight_51_9;
wire signed[31:0]    reg_psum_51_9;
wire signed[31:0]    reg_weight_51_10;
wire signed[31:0]    reg_psum_51_10;
wire signed[31:0]    reg_weight_51_11;
wire signed[31:0]    reg_psum_51_11;
wire signed[31:0]    reg_weight_51_12;
wire signed[31:0]    reg_psum_51_12;
wire signed[31:0]    reg_weight_51_13;
wire signed[31:0]    reg_psum_51_13;
wire signed[31:0]    reg_weight_51_14;
wire signed[31:0]    reg_psum_51_14;
wire signed[31:0]    reg_weight_51_15;
wire signed[31:0]    reg_psum_51_15;
wire signed[31:0]    reg_weight_51_16;
wire signed[31:0]    reg_psum_51_16;
wire signed[31:0]    reg_weight_51_17;
wire signed[31:0]    reg_psum_51_17;
wire signed[31:0]    reg_weight_51_18;
wire signed[31:0]    reg_psum_51_18;
wire signed[31:0]    reg_weight_51_19;
wire signed[31:0]    reg_psum_51_19;
wire signed[31:0]    reg_weight_51_20;
wire signed[31:0]    reg_psum_51_20;
wire signed[31:0]    reg_weight_51_21;
wire signed[31:0]    reg_psum_51_21;
wire signed[31:0]    reg_weight_51_22;
wire signed[31:0]    reg_psum_51_22;
wire signed[31:0]    reg_weight_51_23;
wire signed[31:0]    reg_psum_51_23;
wire signed[31:0]    reg_weight_51_24;
wire signed[31:0]    reg_psum_51_24;
wire signed[31:0]    reg_weight_51_25;
wire signed[31:0]    reg_psum_51_25;
wire signed[31:0]    reg_weight_51_26;
wire signed[31:0]    reg_psum_51_26;
wire signed[31:0]    reg_weight_51_27;
wire signed[31:0]    reg_psum_51_27;
wire signed[31:0]    reg_weight_51_28;
wire signed[31:0]    reg_psum_51_28;
wire signed[31:0]    reg_weight_51_29;
wire signed[31:0]    reg_psum_51_29;
wire signed[31:0]    reg_weight_51_30;
wire signed[31:0]    reg_psum_51_30;
wire signed[31:0]    reg_weight_51_31;
wire signed[31:0]    reg_psum_51_31;
wire signed[31:0]    reg_weight_51_32;
wire signed[31:0]    reg_psum_51_32;
wire signed[31:0]    reg_weight_51_33;
wire signed[31:0]    reg_psum_51_33;
wire signed[31:0]    reg_weight_51_34;
wire signed[31:0]    reg_psum_51_34;
wire signed[31:0]    reg_weight_51_35;
wire signed[31:0]    reg_psum_51_35;
wire signed[31:0]    reg_weight_51_36;
wire signed[31:0]    reg_psum_51_36;
wire signed[31:0]    reg_weight_51_37;
wire signed[31:0]    reg_psum_51_37;
wire signed[31:0]    reg_weight_51_38;
wire signed[31:0]    reg_psum_51_38;
wire signed[31:0]    reg_weight_51_39;
wire signed[31:0]    reg_psum_51_39;
wire signed[31:0]    reg_weight_51_40;
wire signed[31:0]    reg_psum_51_40;
wire signed[31:0]    reg_weight_51_41;
wire signed[31:0]    reg_psum_51_41;
wire signed[31:0]    reg_weight_51_42;
wire signed[31:0]    reg_psum_51_42;
wire signed[31:0]    reg_weight_51_43;
wire signed[31:0]    reg_psum_51_43;
wire signed[31:0]    reg_weight_51_44;
wire signed[31:0]    reg_psum_51_44;
wire signed[31:0]    reg_weight_51_45;
wire signed[31:0]    reg_psum_51_45;
wire signed[31:0]    reg_weight_51_46;
wire signed[31:0]    reg_psum_51_46;
wire signed[31:0]    reg_weight_51_47;
wire signed[31:0]    reg_psum_51_47;
wire signed[31:0]    reg_weight_51_48;
wire signed[31:0]    reg_psum_51_48;
wire signed[31:0]    reg_weight_51_49;
wire signed[31:0]    reg_psum_51_49;
wire signed[31:0]    reg_weight_51_50;
wire signed[31:0]    reg_psum_51_50;
wire signed[31:0]    reg_weight_51_51;
wire signed[31:0]    reg_psum_51_51;
wire signed[31:0]    reg_weight_51_52;
wire signed[31:0]    reg_psum_51_52;
wire signed[31:0]    reg_weight_51_53;
wire signed[31:0]    reg_psum_51_53;
wire signed[31:0]    reg_weight_51_54;
wire signed[31:0]    reg_psum_51_54;
wire signed[31:0]    reg_weight_51_55;
wire signed[31:0]    reg_psum_51_55;
wire signed[31:0]    reg_weight_51_56;
wire signed[31:0]    reg_psum_51_56;
wire signed[31:0]    reg_weight_51_57;
wire signed[31:0]    reg_psum_51_57;
wire signed[31:0]    reg_weight_51_58;
wire signed[31:0]    reg_psum_51_58;
wire signed[31:0]    reg_weight_51_59;
wire signed[31:0]    reg_psum_51_59;
wire signed[31:0]    reg_weight_51_60;
wire signed[31:0]    reg_psum_51_60;
wire signed[31:0]    reg_weight_51_61;
wire signed[31:0]    reg_psum_51_61;
wire signed[31:0]    reg_weight_51_62;
wire signed[31:0]    reg_psum_51_62;
wire signed[31:0]    reg_weight_51_63;
wire signed[31:0]    reg_psum_51_63;
wire signed[31:0]    reg_weight_52_0;
wire signed[31:0]    reg_psum_52_0;
wire signed[31:0]    reg_weight_52_1;
wire signed[31:0]    reg_psum_52_1;
wire signed[31:0]    reg_weight_52_2;
wire signed[31:0]    reg_psum_52_2;
wire signed[31:0]    reg_weight_52_3;
wire signed[31:0]    reg_psum_52_3;
wire signed[31:0]    reg_weight_52_4;
wire signed[31:0]    reg_psum_52_4;
wire signed[31:0]    reg_weight_52_5;
wire signed[31:0]    reg_psum_52_5;
wire signed[31:0]    reg_weight_52_6;
wire signed[31:0]    reg_psum_52_6;
wire signed[31:0]    reg_weight_52_7;
wire signed[31:0]    reg_psum_52_7;
wire signed[31:0]    reg_weight_52_8;
wire signed[31:0]    reg_psum_52_8;
wire signed[31:0]    reg_weight_52_9;
wire signed[31:0]    reg_psum_52_9;
wire signed[31:0]    reg_weight_52_10;
wire signed[31:0]    reg_psum_52_10;
wire signed[31:0]    reg_weight_52_11;
wire signed[31:0]    reg_psum_52_11;
wire signed[31:0]    reg_weight_52_12;
wire signed[31:0]    reg_psum_52_12;
wire signed[31:0]    reg_weight_52_13;
wire signed[31:0]    reg_psum_52_13;
wire signed[31:0]    reg_weight_52_14;
wire signed[31:0]    reg_psum_52_14;
wire signed[31:0]    reg_weight_52_15;
wire signed[31:0]    reg_psum_52_15;
wire signed[31:0]    reg_weight_52_16;
wire signed[31:0]    reg_psum_52_16;
wire signed[31:0]    reg_weight_52_17;
wire signed[31:0]    reg_psum_52_17;
wire signed[31:0]    reg_weight_52_18;
wire signed[31:0]    reg_psum_52_18;
wire signed[31:0]    reg_weight_52_19;
wire signed[31:0]    reg_psum_52_19;
wire signed[31:0]    reg_weight_52_20;
wire signed[31:0]    reg_psum_52_20;
wire signed[31:0]    reg_weight_52_21;
wire signed[31:0]    reg_psum_52_21;
wire signed[31:0]    reg_weight_52_22;
wire signed[31:0]    reg_psum_52_22;
wire signed[31:0]    reg_weight_52_23;
wire signed[31:0]    reg_psum_52_23;
wire signed[31:0]    reg_weight_52_24;
wire signed[31:0]    reg_psum_52_24;
wire signed[31:0]    reg_weight_52_25;
wire signed[31:0]    reg_psum_52_25;
wire signed[31:0]    reg_weight_52_26;
wire signed[31:0]    reg_psum_52_26;
wire signed[31:0]    reg_weight_52_27;
wire signed[31:0]    reg_psum_52_27;
wire signed[31:0]    reg_weight_52_28;
wire signed[31:0]    reg_psum_52_28;
wire signed[31:0]    reg_weight_52_29;
wire signed[31:0]    reg_psum_52_29;
wire signed[31:0]    reg_weight_52_30;
wire signed[31:0]    reg_psum_52_30;
wire signed[31:0]    reg_weight_52_31;
wire signed[31:0]    reg_psum_52_31;
wire signed[31:0]    reg_weight_52_32;
wire signed[31:0]    reg_psum_52_32;
wire signed[31:0]    reg_weight_52_33;
wire signed[31:0]    reg_psum_52_33;
wire signed[31:0]    reg_weight_52_34;
wire signed[31:0]    reg_psum_52_34;
wire signed[31:0]    reg_weight_52_35;
wire signed[31:0]    reg_psum_52_35;
wire signed[31:0]    reg_weight_52_36;
wire signed[31:0]    reg_psum_52_36;
wire signed[31:0]    reg_weight_52_37;
wire signed[31:0]    reg_psum_52_37;
wire signed[31:0]    reg_weight_52_38;
wire signed[31:0]    reg_psum_52_38;
wire signed[31:0]    reg_weight_52_39;
wire signed[31:0]    reg_psum_52_39;
wire signed[31:0]    reg_weight_52_40;
wire signed[31:0]    reg_psum_52_40;
wire signed[31:0]    reg_weight_52_41;
wire signed[31:0]    reg_psum_52_41;
wire signed[31:0]    reg_weight_52_42;
wire signed[31:0]    reg_psum_52_42;
wire signed[31:0]    reg_weight_52_43;
wire signed[31:0]    reg_psum_52_43;
wire signed[31:0]    reg_weight_52_44;
wire signed[31:0]    reg_psum_52_44;
wire signed[31:0]    reg_weight_52_45;
wire signed[31:0]    reg_psum_52_45;
wire signed[31:0]    reg_weight_52_46;
wire signed[31:0]    reg_psum_52_46;
wire signed[31:0]    reg_weight_52_47;
wire signed[31:0]    reg_psum_52_47;
wire signed[31:0]    reg_weight_52_48;
wire signed[31:0]    reg_psum_52_48;
wire signed[31:0]    reg_weight_52_49;
wire signed[31:0]    reg_psum_52_49;
wire signed[31:0]    reg_weight_52_50;
wire signed[31:0]    reg_psum_52_50;
wire signed[31:0]    reg_weight_52_51;
wire signed[31:0]    reg_psum_52_51;
wire signed[31:0]    reg_weight_52_52;
wire signed[31:0]    reg_psum_52_52;
wire signed[31:0]    reg_weight_52_53;
wire signed[31:0]    reg_psum_52_53;
wire signed[31:0]    reg_weight_52_54;
wire signed[31:0]    reg_psum_52_54;
wire signed[31:0]    reg_weight_52_55;
wire signed[31:0]    reg_psum_52_55;
wire signed[31:0]    reg_weight_52_56;
wire signed[31:0]    reg_psum_52_56;
wire signed[31:0]    reg_weight_52_57;
wire signed[31:0]    reg_psum_52_57;
wire signed[31:0]    reg_weight_52_58;
wire signed[31:0]    reg_psum_52_58;
wire signed[31:0]    reg_weight_52_59;
wire signed[31:0]    reg_psum_52_59;
wire signed[31:0]    reg_weight_52_60;
wire signed[31:0]    reg_psum_52_60;
wire signed[31:0]    reg_weight_52_61;
wire signed[31:0]    reg_psum_52_61;
wire signed[31:0]    reg_weight_52_62;
wire signed[31:0]    reg_psum_52_62;
wire signed[31:0]    reg_weight_52_63;
wire signed[31:0]    reg_psum_52_63;
wire signed[31:0]    reg_weight_53_0;
wire signed[31:0]    reg_psum_53_0;
wire signed[31:0]    reg_weight_53_1;
wire signed[31:0]    reg_psum_53_1;
wire signed[31:0]    reg_weight_53_2;
wire signed[31:0]    reg_psum_53_2;
wire signed[31:0]    reg_weight_53_3;
wire signed[31:0]    reg_psum_53_3;
wire signed[31:0]    reg_weight_53_4;
wire signed[31:0]    reg_psum_53_4;
wire signed[31:0]    reg_weight_53_5;
wire signed[31:0]    reg_psum_53_5;
wire signed[31:0]    reg_weight_53_6;
wire signed[31:0]    reg_psum_53_6;
wire signed[31:0]    reg_weight_53_7;
wire signed[31:0]    reg_psum_53_7;
wire signed[31:0]    reg_weight_53_8;
wire signed[31:0]    reg_psum_53_8;
wire signed[31:0]    reg_weight_53_9;
wire signed[31:0]    reg_psum_53_9;
wire signed[31:0]    reg_weight_53_10;
wire signed[31:0]    reg_psum_53_10;
wire signed[31:0]    reg_weight_53_11;
wire signed[31:0]    reg_psum_53_11;
wire signed[31:0]    reg_weight_53_12;
wire signed[31:0]    reg_psum_53_12;
wire signed[31:0]    reg_weight_53_13;
wire signed[31:0]    reg_psum_53_13;
wire signed[31:0]    reg_weight_53_14;
wire signed[31:0]    reg_psum_53_14;
wire signed[31:0]    reg_weight_53_15;
wire signed[31:0]    reg_psum_53_15;
wire signed[31:0]    reg_weight_53_16;
wire signed[31:0]    reg_psum_53_16;
wire signed[31:0]    reg_weight_53_17;
wire signed[31:0]    reg_psum_53_17;
wire signed[31:0]    reg_weight_53_18;
wire signed[31:0]    reg_psum_53_18;
wire signed[31:0]    reg_weight_53_19;
wire signed[31:0]    reg_psum_53_19;
wire signed[31:0]    reg_weight_53_20;
wire signed[31:0]    reg_psum_53_20;
wire signed[31:0]    reg_weight_53_21;
wire signed[31:0]    reg_psum_53_21;
wire signed[31:0]    reg_weight_53_22;
wire signed[31:0]    reg_psum_53_22;
wire signed[31:0]    reg_weight_53_23;
wire signed[31:0]    reg_psum_53_23;
wire signed[31:0]    reg_weight_53_24;
wire signed[31:0]    reg_psum_53_24;
wire signed[31:0]    reg_weight_53_25;
wire signed[31:0]    reg_psum_53_25;
wire signed[31:0]    reg_weight_53_26;
wire signed[31:0]    reg_psum_53_26;
wire signed[31:0]    reg_weight_53_27;
wire signed[31:0]    reg_psum_53_27;
wire signed[31:0]    reg_weight_53_28;
wire signed[31:0]    reg_psum_53_28;
wire signed[31:0]    reg_weight_53_29;
wire signed[31:0]    reg_psum_53_29;
wire signed[31:0]    reg_weight_53_30;
wire signed[31:0]    reg_psum_53_30;
wire signed[31:0]    reg_weight_53_31;
wire signed[31:0]    reg_psum_53_31;
wire signed[31:0]    reg_weight_53_32;
wire signed[31:0]    reg_psum_53_32;
wire signed[31:0]    reg_weight_53_33;
wire signed[31:0]    reg_psum_53_33;
wire signed[31:0]    reg_weight_53_34;
wire signed[31:0]    reg_psum_53_34;
wire signed[31:0]    reg_weight_53_35;
wire signed[31:0]    reg_psum_53_35;
wire signed[31:0]    reg_weight_53_36;
wire signed[31:0]    reg_psum_53_36;
wire signed[31:0]    reg_weight_53_37;
wire signed[31:0]    reg_psum_53_37;
wire signed[31:0]    reg_weight_53_38;
wire signed[31:0]    reg_psum_53_38;
wire signed[31:0]    reg_weight_53_39;
wire signed[31:0]    reg_psum_53_39;
wire signed[31:0]    reg_weight_53_40;
wire signed[31:0]    reg_psum_53_40;
wire signed[31:0]    reg_weight_53_41;
wire signed[31:0]    reg_psum_53_41;
wire signed[31:0]    reg_weight_53_42;
wire signed[31:0]    reg_psum_53_42;
wire signed[31:0]    reg_weight_53_43;
wire signed[31:0]    reg_psum_53_43;
wire signed[31:0]    reg_weight_53_44;
wire signed[31:0]    reg_psum_53_44;
wire signed[31:0]    reg_weight_53_45;
wire signed[31:0]    reg_psum_53_45;
wire signed[31:0]    reg_weight_53_46;
wire signed[31:0]    reg_psum_53_46;
wire signed[31:0]    reg_weight_53_47;
wire signed[31:0]    reg_psum_53_47;
wire signed[31:0]    reg_weight_53_48;
wire signed[31:0]    reg_psum_53_48;
wire signed[31:0]    reg_weight_53_49;
wire signed[31:0]    reg_psum_53_49;
wire signed[31:0]    reg_weight_53_50;
wire signed[31:0]    reg_psum_53_50;
wire signed[31:0]    reg_weight_53_51;
wire signed[31:0]    reg_psum_53_51;
wire signed[31:0]    reg_weight_53_52;
wire signed[31:0]    reg_psum_53_52;
wire signed[31:0]    reg_weight_53_53;
wire signed[31:0]    reg_psum_53_53;
wire signed[31:0]    reg_weight_53_54;
wire signed[31:0]    reg_psum_53_54;
wire signed[31:0]    reg_weight_53_55;
wire signed[31:0]    reg_psum_53_55;
wire signed[31:0]    reg_weight_53_56;
wire signed[31:0]    reg_psum_53_56;
wire signed[31:0]    reg_weight_53_57;
wire signed[31:0]    reg_psum_53_57;
wire signed[31:0]    reg_weight_53_58;
wire signed[31:0]    reg_psum_53_58;
wire signed[31:0]    reg_weight_53_59;
wire signed[31:0]    reg_psum_53_59;
wire signed[31:0]    reg_weight_53_60;
wire signed[31:0]    reg_psum_53_60;
wire signed[31:0]    reg_weight_53_61;
wire signed[31:0]    reg_psum_53_61;
wire signed[31:0]    reg_weight_53_62;
wire signed[31:0]    reg_psum_53_62;
wire signed[31:0]    reg_weight_53_63;
wire signed[31:0]    reg_psum_53_63;
wire signed[31:0]    reg_weight_54_0;
wire signed[31:0]    reg_psum_54_0;
wire signed[31:0]    reg_weight_54_1;
wire signed[31:0]    reg_psum_54_1;
wire signed[31:0]    reg_weight_54_2;
wire signed[31:0]    reg_psum_54_2;
wire signed[31:0]    reg_weight_54_3;
wire signed[31:0]    reg_psum_54_3;
wire signed[31:0]    reg_weight_54_4;
wire signed[31:0]    reg_psum_54_4;
wire signed[31:0]    reg_weight_54_5;
wire signed[31:0]    reg_psum_54_5;
wire signed[31:0]    reg_weight_54_6;
wire signed[31:0]    reg_psum_54_6;
wire signed[31:0]    reg_weight_54_7;
wire signed[31:0]    reg_psum_54_7;
wire signed[31:0]    reg_weight_54_8;
wire signed[31:0]    reg_psum_54_8;
wire signed[31:0]    reg_weight_54_9;
wire signed[31:0]    reg_psum_54_9;
wire signed[31:0]    reg_weight_54_10;
wire signed[31:0]    reg_psum_54_10;
wire signed[31:0]    reg_weight_54_11;
wire signed[31:0]    reg_psum_54_11;
wire signed[31:0]    reg_weight_54_12;
wire signed[31:0]    reg_psum_54_12;
wire signed[31:0]    reg_weight_54_13;
wire signed[31:0]    reg_psum_54_13;
wire signed[31:0]    reg_weight_54_14;
wire signed[31:0]    reg_psum_54_14;
wire signed[31:0]    reg_weight_54_15;
wire signed[31:0]    reg_psum_54_15;
wire signed[31:0]    reg_weight_54_16;
wire signed[31:0]    reg_psum_54_16;
wire signed[31:0]    reg_weight_54_17;
wire signed[31:0]    reg_psum_54_17;
wire signed[31:0]    reg_weight_54_18;
wire signed[31:0]    reg_psum_54_18;
wire signed[31:0]    reg_weight_54_19;
wire signed[31:0]    reg_psum_54_19;
wire signed[31:0]    reg_weight_54_20;
wire signed[31:0]    reg_psum_54_20;
wire signed[31:0]    reg_weight_54_21;
wire signed[31:0]    reg_psum_54_21;
wire signed[31:0]    reg_weight_54_22;
wire signed[31:0]    reg_psum_54_22;
wire signed[31:0]    reg_weight_54_23;
wire signed[31:0]    reg_psum_54_23;
wire signed[31:0]    reg_weight_54_24;
wire signed[31:0]    reg_psum_54_24;
wire signed[31:0]    reg_weight_54_25;
wire signed[31:0]    reg_psum_54_25;
wire signed[31:0]    reg_weight_54_26;
wire signed[31:0]    reg_psum_54_26;
wire signed[31:0]    reg_weight_54_27;
wire signed[31:0]    reg_psum_54_27;
wire signed[31:0]    reg_weight_54_28;
wire signed[31:0]    reg_psum_54_28;
wire signed[31:0]    reg_weight_54_29;
wire signed[31:0]    reg_psum_54_29;
wire signed[31:0]    reg_weight_54_30;
wire signed[31:0]    reg_psum_54_30;
wire signed[31:0]    reg_weight_54_31;
wire signed[31:0]    reg_psum_54_31;
wire signed[31:0]    reg_weight_54_32;
wire signed[31:0]    reg_psum_54_32;
wire signed[31:0]    reg_weight_54_33;
wire signed[31:0]    reg_psum_54_33;
wire signed[31:0]    reg_weight_54_34;
wire signed[31:0]    reg_psum_54_34;
wire signed[31:0]    reg_weight_54_35;
wire signed[31:0]    reg_psum_54_35;
wire signed[31:0]    reg_weight_54_36;
wire signed[31:0]    reg_psum_54_36;
wire signed[31:0]    reg_weight_54_37;
wire signed[31:0]    reg_psum_54_37;
wire signed[31:0]    reg_weight_54_38;
wire signed[31:0]    reg_psum_54_38;
wire signed[31:0]    reg_weight_54_39;
wire signed[31:0]    reg_psum_54_39;
wire signed[31:0]    reg_weight_54_40;
wire signed[31:0]    reg_psum_54_40;
wire signed[31:0]    reg_weight_54_41;
wire signed[31:0]    reg_psum_54_41;
wire signed[31:0]    reg_weight_54_42;
wire signed[31:0]    reg_psum_54_42;
wire signed[31:0]    reg_weight_54_43;
wire signed[31:0]    reg_psum_54_43;
wire signed[31:0]    reg_weight_54_44;
wire signed[31:0]    reg_psum_54_44;
wire signed[31:0]    reg_weight_54_45;
wire signed[31:0]    reg_psum_54_45;
wire signed[31:0]    reg_weight_54_46;
wire signed[31:0]    reg_psum_54_46;
wire signed[31:0]    reg_weight_54_47;
wire signed[31:0]    reg_psum_54_47;
wire signed[31:0]    reg_weight_54_48;
wire signed[31:0]    reg_psum_54_48;
wire signed[31:0]    reg_weight_54_49;
wire signed[31:0]    reg_psum_54_49;
wire signed[31:0]    reg_weight_54_50;
wire signed[31:0]    reg_psum_54_50;
wire signed[31:0]    reg_weight_54_51;
wire signed[31:0]    reg_psum_54_51;
wire signed[31:0]    reg_weight_54_52;
wire signed[31:0]    reg_psum_54_52;
wire signed[31:0]    reg_weight_54_53;
wire signed[31:0]    reg_psum_54_53;
wire signed[31:0]    reg_weight_54_54;
wire signed[31:0]    reg_psum_54_54;
wire signed[31:0]    reg_weight_54_55;
wire signed[31:0]    reg_psum_54_55;
wire signed[31:0]    reg_weight_54_56;
wire signed[31:0]    reg_psum_54_56;
wire signed[31:0]    reg_weight_54_57;
wire signed[31:0]    reg_psum_54_57;
wire signed[31:0]    reg_weight_54_58;
wire signed[31:0]    reg_psum_54_58;
wire signed[31:0]    reg_weight_54_59;
wire signed[31:0]    reg_psum_54_59;
wire signed[31:0]    reg_weight_54_60;
wire signed[31:0]    reg_psum_54_60;
wire signed[31:0]    reg_weight_54_61;
wire signed[31:0]    reg_psum_54_61;
wire signed[31:0]    reg_weight_54_62;
wire signed[31:0]    reg_psum_54_62;
wire signed[31:0]    reg_weight_54_63;
wire signed[31:0]    reg_psum_54_63;
wire signed[31:0]    reg_weight_55_0;
wire signed[31:0]    reg_psum_55_0;
wire signed[31:0]    reg_weight_55_1;
wire signed[31:0]    reg_psum_55_1;
wire signed[31:0]    reg_weight_55_2;
wire signed[31:0]    reg_psum_55_2;
wire signed[31:0]    reg_weight_55_3;
wire signed[31:0]    reg_psum_55_3;
wire signed[31:0]    reg_weight_55_4;
wire signed[31:0]    reg_psum_55_4;
wire signed[31:0]    reg_weight_55_5;
wire signed[31:0]    reg_psum_55_5;
wire signed[31:0]    reg_weight_55_6;
wire signed[31:0]    reg_psum_55_6;
wire signed[31:0]    reg_weight_55_7;
wire signed[31:0]    reg_psum_55_7;
wire signed[31:0]    reg_weight_55_8;
wire signed[31:0]    reg_psum_55_8;
wire signed[31:0]    reg_weight_55_9;
wire signed[31:0]    reg_psum_55_9;
wire signed[31:0]    reg_weight_55_10;
wire signed[31:0]    reg_psum_55_10;
wire signed[31:0]    reg_weight_55_11;
wire signed[31:0]    reg_psum_55_11;
wire signed[31:0]    reg_weight_55_12;
wire signed[31:0]    reg_psum_55_12;
wire signed[31:0]    reg_weight_55_13;
wire signed[31:0]    reg_psum_55_13;
wire signed[31:0]    reg_weight_55_14;
wire signed[31:0]    reg_psum_55_14;
wire signed[31:0]    reg_weight_55_15;
wire signed[31:0]    reg_psum_55_15;
wire signed[31:0]    reg_weight_55_16;
wire signed[31:0]    reg_psum_55_16;
wire signed[31:0]    reg_weight_55_17;
wire signed[31:0]    reg_psum_55_17;
wire signed[31:0]    reg_weight_55_18;
wire signed[31:0]    reg_psum_55_18;
wire signed[31:0]    reg_weight_55_19;
wire signed[31:0]    reg_psum_55_19;
wire signed[31:0]    reg_weight_55_20;
wire signed[31:0]    reg_psum_55_20;
wire signed[31:0]    reg_weight_55_21;
wire signed[31:0]    reg_psum_55_21;
wire signed[31:0]    reg_weight_55_22;
wire signed[31:0]    reg_psum_55_22;
wire signed[31:0]    reg_weight_55_23;
wire signed[31:0]    reg_psum_55_23;
wire signed[31:0]    reg_weight_55_24;
wire signed[31:0]    reg_psum_55_24;
wire signed[31:0]    reg_weight_55_25;
wire signed[31:0]    reg_psum_55_25;
wire signed[31:0]    reg_weight_55_26;
wire signed[31:0]    reg_psum_55_26;
wire signed[31:0]    reg_weight_55_27;
wire signed[31:0]    reg_psum_55_27;
wire signed[31:0]    reg_weight_55_28;
wire signed[31:0]    reg_psum_55_28;
wire signed[31:0]    reg_weight_55_29;
wire signed[31:0]    reg_psum_55_29;
wire signed[31:0]    reg_weight_55_30;
wire signed[31:0]    reg_psum_55_30;
wire signed[31:0]    reg_weight_55_31;
wire signed[31:0]    reg_psum_55_31;
wire signed[31:0]    reg_weight_55_32;
wire signed[31:0]    reg_psum_55_32;
wire signed[31:0]    reg_weight_55_33;
wire signed[31:0]    reg_psum_55_33;
wire signed[31:0]    reg_weight_55_34;
wire signed[31:0]    reg_psum_55_34;
wire signed[31:0]    reg_weight_55_35;
wire signed[31:0]    reg_psum_55_35;
wire signed[31:0]    reg_weight_55_36;
wire signed[31:0]    reg_psum_55_36;
wire signed[31:0]    reg_weight_55_37;
wire signed[31:0]    reg_psum_55_37;
wire signed[31:0]    reg_weight_55_38;
wire signed[31:0]    reg_psum_55_38;
wire signed[31:0]    reg_weight_55_39;
wire signed[31:0]    reg_psum_55_39;
wire signed[31:0]    reg_weight_55_40;
wire signed[31:0]    reg_psum_55_40;
wire signed[31:0]    reg_weight_55_41;
wire signed[31:0]    reg_psum_55_41;
wire signed[31:0]    reg_weight_55_42;
wire signed[31:0]    reg_psum_55_42;
wire signed[31:0]    reg_weight_55_43;
wire signed[31:0]    reg_psum_55_43;
wire signed[31:0]    reg_weight_55_44;
wire signed[31:0]    reg_psum_55_44;
wire signed[31:0]    reg_weight_55_45;
wire signed[31:0]    reg_psum_55_45;
wire signed[31:0]    reg_weight_55_46;
wire signed[31:0]    reg_psum_55_46;
wire signed[31:0]    reg_weight_55_47;
wire signed[31:0]    reg_psum_55_47;
wire signed[31:0]    reg_weight_55_48;
wire signed[31:0]    reg_psum_55_48;
wire signed[31:0]    reg_weight_55_49;
wire signed[31:0]    reg_psum_55_49;
wire signed[31:0]    reg_weight_55_50;
wire signed[31:0]    reg_psum_55_50;
wire signed[31:0]    reg_weight_55_51;
wire signed[31:0]    reg_psum_55_51;
wire signed[31:0]    reg_weight_55_52;
wire signed[31:0]    reg_psum_55_52;
wire signed[31:0]    reg_weight_55_53;
wire signed[31:0]    reg_psum_55_53;
wire signed[31:0]    reg_weight_55_54;
wire signed[31:0]    reg_psum_55_54;
wire signed[31:0]    reg_weight_55_55;
wire signed[31:0]    reg_psum_55_55;
wire signed[31:0]    reg_weight_55_56;
wire signed[31:0]    reg_psum_55_56;
wire signed[31:0]    reg_weight_55_57;
wire signed[31:0]    reg_psum_55_57;
wire signed[31:0]    reg_weight_55_58;
wire signed[31:0]    reg_psum_55_58;
wire signed[31:0]    reg_weight_55_59;
wire signed[31:0]    reg_psum_55_59;
wire signed[31:0]    reg_weight_55_60;
wire signed[31:0]    reg_psum_55_60;
wire signed[31:0]    reg_weight_55_61;
wire signed[31:0]    reg_psum_55_61;
wire signed[31:0]    reg_weight_55_62;
wire signed[31:0]    reg_psum_55_62;
wire signed[31:0]    reg_weight_55_63;
wire signed[31:0]    reg_psum_55_63;
wire signed[31:0]    reg_weight_56_0;
wire signed[31:0]    reg_psum_56_0;
wire signed[31:0]    reg_weight_56_1;
wire signed[31:0]    reg_psum_56_1;
wire signed[31:0]    reg_weight_56_2;
wire signed[31:0]    reg_psum_56_2;
wire signed[31:0]    reg_weight_56_3;
wire signed[31:0]    reg_psum_56_3;
wire signed[31:0]    reg_weight_56_4;
wire signed[31:0]    reg_psum_56_4;
wire signed[31:0]    reg_weight_56_5;
wire signed[31:0]    reg_psum_56_5;
wire signed[31:0]    reg_weight_56_6;
wire signed[31:0]    reg_psum_56_6;
wire signed[31:0]    reg_weight_56_7;
wire signed[31:0]    reg_psum_56_7;
wire signed[31:0]    reg_weight_56_8;
wire signed[31:0]    reg_psum_56_8;
wire signed[31:0]    reg_weight_56_9;
wire signed[31:0]    reg_psum_56_9;
wire signed[31:0]    reg_weight_56_10;
wire signed[31:0]    reg_psum_56_10;
wire signed[31:0]    reg_weight_56_11;
wire signed[31:0]    reg_psum_56_11;
wire signed[31:0]    reg_weight_56_12;
wire signed[31:0]    reg_psum_56_12;
wire signed[31:0]    reg_weight_56_13;
wire signed[31:0]    reg_psum_56_13;
wire signed[31:0]    reg_weight_56_14;
wire signed[31:0]    reg_psum_56_14;
wire signed[31:0]    reg_weight_56_15;
wire signed[31:0]    reg_psum_56_15;
wire signed[31:0]    reg_weight_56_16;
wire signed[31:0]    reg_psum_56_16;
wire signed[31:0]    reg_weight_56_17;
wire signed[31:0]    reg_psum_56_17;
wire signed[31:0]    reg_weight_56_18;
wire signed[31:0]    reg_psum_56_18;
wire signed[31:0]    reg_weight_56_19;
wire signed[31:0]    reg_psum_56_19;
wire signed[31:0]    reg_weight_56_20;
wire signed[31:0]    reg_psum_56_20;
wire signed[31:0]    reg_weight_56_21;
wire signed[31:0]    reg_psum_56_21;
wire signed[31:0]    reg_weight_56_22;
wire signed[31:0]    reg_psum_56_22;
wire signed[31:0]    reg_weight_56_23;
wire signed[31:0]    reg_psum_56_23;
wire signed[31:0]    reg_weight_56_24;
wire signed[31:0]    reg_psum_56_24;
wire signed[31:0]    reg_weight_56_25;
wire signed[31:0]    reg_psum_56_25;
wire signed[31:0]    reg_weight_56_26;
wire signed[31:0]    reg_psum_56_26;
wire signed[31:0]    reg_weight_56_27;
wire signed[31:0]    reg_psum_56_27;
wire signed[31:0]    reg_weight_56_28;
wire signed[31:0]    reg_psum_56_28;
wire signed[31:0]    reg_weight_56_29;
wire signed[31:0]    reg_psum_56_29;
wire signed[31:0]    reg_weight_56_30;
wire signed[31:0]    reg_psum_56_30;
wire signed[31:0]    reg_weight_56_31;
wire signed[31:0]    reg_psum_56_31;
wire signed[31:0]    reg_weight_56_32;
wire signed[31:0]    reg_psum_56_32;
wire signed[31:0]    reg_weight_56_33;
wire signed[31:0]    reg_psum_56_33;
wire signed[31:0]    reg_weight_56_34;
wire signed[31:0]    reg_psum_56_34;
wire signed[31:0]    reg_weight_56_35;
wire signed[31:0]    reg_psum_56_35;
wire signed[31:0]    reg_weight_56_36;
wire signed[31:0]    reg_psum_56_36;
wire signed[31:0]    reg_weight_56_37;
wire signed[31:0]    reg_psum_56_37;
wire signed[31:0]    reg_weight_56_38;
wire signed[31:0]    reg_psum_56_38;
wire signed[31:0]    reg_weight_56_39;
wire signed[31:0]    reg_psum_56_39;
wire signed[31:0]    reg_weight_56_40;
wire signed[31:0]    reg_psum_56_40;
wire signed[31:0]    reg_weight_56_41;
wire signed[31:0]    reg_psum_56_41;
wire signed[31:0]    reg_weight_56_42;
wire signed[31:0]    reg_psum_56_42;
wire signed[31:0]    reg_weight_56_43;
wire signed[31:0]    reg_psum_56_43;
wire signed[31:0]    reg_weight_56_44;
wire signed[31:0]    reg_psum_56_44;
wire signed[31:0]    reg_weight_56_45;
wire signed[31:0]    reg_psum_56_45;
wire signed[31:0]    reg_weight_56_46;
wire signed[31:0]    reg_psum_56_46;
wire signed[31:0]    reg_weight_56_47;
wire signed[31:0]    reg_psum_56_47;
wire signed[31:0]    reg_weight_56_48;
wire signed[31:0]    reg_psum_56_48;
wire signed[31:0]    reg_weight_56_49;
wire signed[31:0]    reg_psum_56_49;
wire signed[31:0]    reg_weight_56_50;
wire signed[31:0]    reg_psum_56_50;
wire signed[31:0]    reg_weight_56_51;
wire signed[31:0]    reg_psum_56_51;
wire signed[31:0]    reg_weight_56_52;
wire signed[31:0]    reg_psum_56_52;
wire signed[31:0]    reg_weight_56_53;
wire signed[31:0]    reg_psum_56_53;
wire signed[31:0]    reg_weight_56_54;
wire signed[31:0]    reg_psum_56_54;
wire signed[31:0]    reg_weight_56_55;
wire signed[31:0]    reg_psum_56_55;
wire signed[31:0]    reg_weight_56_56;
wire signed[31:0]    reg_psum_56_56;
wire signed[31:0]    reg_weight_56_57;
wire signed[31:0]    reg_psum_56_57;
wire signed[31:0]    reg_weight_56_58;
wire signed[31:0]    reg_psum_56_58;
wire signed[31:0]    reg_weight_56_59;
wire signed[31:0]    reg_psum_56_59;
wire signed[31:0]    reg_weight_56_60;
wire signed[31:0]    reg_psum_56_60;
wire signed[31:0]    reg_weight_56_61;
wire signed[31:0]    reg_psum_56_61;
wire signed[31:0]    reg_weight_56_62;
wire signed[31:0]    reg_psum_56_62;
wire signed[31:0]    reg_weight_56_63;
wire signed[31:0]    reg_psum_56_63;
wire signed[31:0]    reg_weight_57_0;
wire signed[31:0]    reg_psum_57_0;
wire signed[31:0]    reg_weight_57_1;
wire signed[31:0]    reg_psum_57_1;
wire signed[31:0]    reg_weight_57_2;
wire signed[31:0]    reg_psum_57_2;
wire signed[31:0]    reg_weight_57_3;
wire signed[31:0]    reg_psum_57_3;
wire signed[31:0]    reg_weight_57_4;
wire signed[31:0]    reg_psum_57_4;
wire signed[31:0]    reg_weight_57_5;
wire signed[31:0]    reg_psum_57_5;
wire signed[31:0]    reg_weight_57_6;
wire signed[31:0]    reg_psum_57_6;
wire signed[31:0]    reg_weight_57_7;
wire signed[31:0]    reg_psum_57_7;
wire signed[31:0]    reg_weight_57_8;
wire signed[31:0]    reg_psum_57_8;
wire signed[31:0]    reg_weight_57_9;
wire signed[31:0]    reg_psum_57_9;
wire signed[31:0]    reg_weight_57_10;
wire signed[31:0]    reg_psum_57_10;
wire signed[31:0]    reg_weight_57_11;
wire signed[31:0]    reg_psum_57_11;
wire signed[31:0]    reg_weight_57_12;
wire signed[31:0]    reg_psum_57_12;
wire signed[31:0]    reg_weight_57_13;
wire signed[31:0]    reg_psum_57_13;
wire signed[31:0]    reg_weight_57_14;
wire signed[31:0]    reg_psum_57_14;
wire signed[31:0]    reg_weight_57_15;
wire signed[31:0]    reg_psum_57_15;
wire signed[31:0]    reg_weight_57_16;
wire signed[31:0]    reg_psum_57_16;
wire signed[31:0]    reg_weight_57_17;
wire signed[31:0]    reg_psum_57_17;
wire signed[31:0]    reg_weight_57_18;
wire signed[31:0]    reg_psum_57_18;
wire signed[31:0]    reg_weight_57_19;
wire signed[31:0]    reg_psum_57_19;
wire signed[31:0]    reg_weight_57_20;
wire signed[31:0]    reg_psum_57_20;
wire signed[31:0]    reg_weight_57_21;
wire signed[31:0]    reg_psum_57_21;
wire signed[31:0]    reg_weight_57_22;
wire signed[31:0]    reg_psum_57_22;
wire signed[31:0]    reg_weight_57_23;
wire signed[31:0]    reg_psum_57_23;
wire signed[31:0]    reg_weight_57_24;
wire signed[31:0]    reg_psum_57_24;
wire signed[31:0]    reg_weight_57_25;
wire signed[31:0]    reg_psum_57_25;
wire signed[31:0]    reg_weight_57_26;
wire signed[31:0]    reg_psum_57_26;
wire signed[31:0]    reg_weight_57_27;
wire signed[31:0]    reg_psum_57_27;
wire signed[31:0]    reg_weight_57_28;
wire signed[31:0]    reg_psum_57_28;
wire signed[31:0]    reg_weight_57_29;
wire signed[31:0]    reg_psum_57_29;
wire signed[31:0]    reg_weight_57_30;
wire signed[31:0]    reg_psum_57_30;
wire signed[31:0]    reg_weight_57_31;
wire signed[31:0]    reg_psum_57_31;
wire signed[31:0]    reg_weight_57_32;
wire signed[31:0]    reg_psum_57_32;
wire signed[31:0]    reg_weight_57_33;
wire signed[31:0]    reg_psum_57_33;
wire signed[31:0]    reg_weight_57_34;
wire signed[31:0]    reg_psum_57_34;
wire signed[31:0]    reg_weight_57_35;
wire signed[31:0]    reg_psum_57_35;
wire signed[31:0]    reg_weight_57_36;
wire signed[31:0]    reg_psum_57_36;
wire signed[31:0]    reg_weight_57_37;
wire signed[31:0]    reg_psum_57_37;
wire signed[31:0]    reg_weight_57_38;
wire signed[31:0]    reg_psum_57_38;
wire signed[31:0]    reg_weight_57_39;
wire signed[31:0]    reg_psum_57_39;
wire signed[31:0]    reg_weight_57_40;
wire signed[31:0]    reg_psum_57_40;
wire signed[31:0]    reg_weight_57_41;
wire signed[31:0]    reg_psum_57_41;
wire signed[31:0]    reg_weight_57_42;
wire signed[31:0]    reg_psum_57_42;
wire signed[31:0]    reg_weight_57_43;
wire signed[31:0]    reg_psum_57_43;
wire signed[31:0]    reg_weight_57_44;
wire signed[31:0]    reg_psum_57_44;
wire signed[31:0]    reg_weight_57_45;
wire signed[31:0]    reg_psum_57_45;
wire signed[31:0]    reg_weight_57_46;
wire signed[31:0]    reg_psum_57_46;
wire signed[31:0]    reg_weight_57_47;
wire signed[31:0]    reg_psum_57_47;
wire signed[31:0]    reg_weight_57_48;
wire signed[31:0]    reg_psum_57_48;
wire signed[31:0]    reg_weight_57_49;
wire signed[31:0]    reg_psum_57_49;
wire signed[31:0]    reg_weight_57_50;
wire signed[31:0]    reg_psum_57_50;
wire signed[31:0]    reg_weight_57_51;
wire signed[31:0]    reg_psum_57_51;
wire signed[31:0]    reg_weight_57_52;
wire signed[31:0]    reg_psum_57_52;
wire signed[31:0]    reg_weight_57_53;
wire signed[31:0]    reg_psum_57_53;
wire signed[31:0]    reg_weight_57_54;
wire signed[31:0]    reg_psum_57_54;
wire signed[31:0]    reg_weight_57_55;
wire signed[31:0]    reg_psum_57_55;
wire signed[31:0]    reg_weight_57_56;
wire signed[31:0]    reg_psum_57_56;
wire signed[31:0]    reg_weight_57_57;
wire signed[31:0]    reg_psum_57_57;
wire signed[31:0]    reg_weight_57_58;
wire signed[31:0]    reg_psum_57_58;
wire signed[31:0]    reg_weight_57_59;
wire signed[31:0]    reg_psum_57_59;
wire signed[31:0]    reg_weight_57_60;
wire signed[31:0]    reg_psum_57_60;
wire signed[31:0]    reg_weight_57_61;
wire signed[31:0]    reg_psum_57_61;
wire signed[31:0]    reg_weight_57_62;
wire signed[31:0]    reg_psum_57_62;
wire signed[31:0]    reg_weight_57_63;
wire signed[31:0]    reg_psum_57_63;
wire signed[31:0]    reg_weight_58_0;
wire signed[31:0]    reg_psum_58_0;
wire signed[31:0]    reg_weight_58_1;
wire signed[31:0]    reg_psum_58_1;
wire signed[31:0]    reg_weight_58_2;
wire signed[31:0]    reg_psum_58_2;
wire signed[31:0]    reg_weight_58_3;
wire signed[31:0]    reg_psum_58_3;
wire signed[31:0]    reg_weight_58_4;
wire signed[31:0]    reg_psum_58_4;
wire signed[31:0]    reg_weight_58_5;
wire signed[31:0]    reg_psum_58_5;
wire signed[31:0]    reg_weight_58_6;
wire signed[31:0]    reg_psum_58_6;
wire signed[31:0]    reg_weight_58_7;
wire signed[31:0]    reg_psum_58_7;
wire signed[31:0]    reg_weight_58_8;
wire signed[31:0]    reg_psum_58_8;
wire signed[31:0]    reg_weight_58_9;
wire signed[31:0]    reg_psum_58_9;
wire signed[31:0]    reg_weight_58_10;
wire signed[31:0]    reg_psum_58_10;
wire signed[31:0]    reg_weight_58_11;
wire signed[31:0]    reg_psum_58_11;
wire signed[31:0]    reg_weight_58_12;
wire signed[31:0]    reg_psum_58_12;
wire signed[31:0]    reg_weight_58_13;
wire signed[31:0]    reg_psum_58_13;
wire signed[31:0]    reg_weight_58_14;
wire signed[31:0]    reg_psum_58_14;
wire signed[31:0]    reg_weight_58_15;
wire signed[31:0]    reg_psum_58_15;
wire signed[31:0]    reg_weight_58_16;
wire signed[31:0]    reg_psum_58_16;
wire signed[31:0]    reg_weight_58_17;
wire signed[31:0]    reg_psum_58_17;
wire signed[31:0]    reg_weight_58_18;
wire signed[31:0]    reg_psum_58_18;
wire signed[31:0]    reg_weight_58_19;
wire signed[31:0]    reg_psum_58_19;
wire signed[31:0]    reg_weight_58_20;
wire signed[31:0]    reg_psum_58_20;
wire signed[31:0]    reg_weight_58_21;
wire signed[31:0]    reg_psum_58_21;
wire signed[31:0]    reg_weight_58_22;
wire signed[31:0]    reg_psum_58_22;
wire signed[31:0]    reg_weight_58_23;
wire signed[31:0]    reg_psum_58_23;
wire signed[31:0]    reg_weight_58_24;
wire signed[31:0]    reg_psum_58_24;
wire signed[31:0]    reg_weight_58_25;
wire signed[31:0]    reg_psum_58_25;
wire signed[31:0]    reg_weight_58_26;
wire signed[31:0]    reg_psum_58_26;
wire signed[31:0]    reg_weight_58_27;
wire signed[31:0]    reg_psum_58_27;
wire signed[31:0]    reg_weight_58_28;
wire signed[31:0]    reg_psum_58_28;
wire signed[31:0]    reg_weight_58_29;
wire signed[31:0]    reg_psum_58_29;
wire signed[31:0]    reg_weight_58_30;
wire signed[31:0]    reg_psum_58_30;
wire signed[31:0]    reg_weight_58_31;
wire signed[31:0]    reg_psum_58_31;
wire signed[31:0]    reg_weight_58_32;
wire signed[31:0]    reg_psum_58_32;
wire signed[31:0]    reg_weight_58_33;
wire signed[31:0]    reg_psum_58_33;
wire signed[31:0]    reg_weight_58_34;
wire signed[31:0]    reg_psum_58_34;
wire signed[31:0]    reg_weight_58_35;
wire signed[31:0]    reg_psum_58_35;
wire signed[31:0]    reg_weight_58_36;
wire signed[31:0]    reg_psum_58_36;
wire signed[31:0]    reg_weight_58_37;
wire signed[31:0]    reg_psum_58_37;
wire signed[31:0]    reg_weight_58_38;
wire signed[31:0]    reg_psum_58_38;
wire signed[31:0]    reg_weight_58_39;
wire signed[31:0]    reg_psum_58_39;
wire signed[31:0]    reg_weight_58_40;
wire signed[31:0]    reg_psum_58_40;
wire signed[31:0]    reg_weight_58_41;
wire signed[31:0]    reg_psum_58_41;
wire signed[31:0]    reg_weight_58_42;
wire signed[31:0]    reg_psum_58_42;
wire signed[31:0]    reg_weight_58_43;
wire signed[31:0]    reg_psum_58_43;
wire signed[31:0]    reg_weight_58_44;
wire signed[31:0]    reg_psum_58_44;
wire signed[31:0]    reg_weight_58_45;
wire signed[31:0]    reg_psum_58_45;
wire signed[31:0]    reg_weight_58_46;
wire signed[31:0]    reg_psum_58_46;
wire signed[31:0]    reg_weight_58_47;
wire signed[31:0]    reg_psum_58_47;
wire signed[31:0]    reg_weight_58_48;
wire signed[31:0]    reg_psum_58_48;
wire signed[31:0]    reg_weight_58_49;
wire signed[31:0]    reg_psum_58_49;
wire signed[31:0]    reg_weight_58_50;
wire signed[31:0]    reg_psum_58_50;
wire signed[31:0]    reg_weight_58_51;
wire signed[31:0]    reg_psum_58_51;
wire signed[31:0]    reg_weight_58_52;
wire signed[31:0]    reg_psum_58_52;
wire signed[31:0]    reg_weight_58_53;
wire signed[31:0]    reg_psum_58_53;
wire signed[31:0]    reg_weight_58_54;
wire signed[31:0]    reg_psum_58_54;
wire signed[31:0]    reg_weight_58_55;
wire signed[31:0]    reg_psum_58_55;
wire signed[31:0]    reg_weight_58_56;
wire signed[31:0]    reg_psum_58_56;
wire signed[31:0]    reg_weight_58_57;
wire signed[31:0]    reg_psum_58_57;
wire signed[31:0]    reg_weight_58_58;
wire signed[31:0]    reg_psum_58_58;
wire signed[31:0]    reg_weight_58_59;
wire signed[31:0]    reg_psum_58_59;
wire signed[31:0]    reg_weight_58_60;
wire signed[31:0]    reg_psum_58_60;
wire signed[31:0]    reg_weight_58_61;
wire signed[31:0]    reg_psum_58_61;
wire signed[31:0]    reg_weight_58_62;
wire signed[31:0]    reg_psum_58_62;
wire signed[31:0]    reg_weight_58_63;
wire signed[31:0]    reg_psum_58_63;
wire signed[31:0]    reg_weight_59_0;
wire signed[31:0]    reg_psum_59_0;
wire signed[31:0]    reg_weight_59_1;
wire signed[31:0]    reg_psum_59_1;
wire signed[31:0]    reg_weight_59_2;
wire signed[31:0]    reg_psum_59_2;
wire signed[31:0]    reg_weight_59_3;
wire signed[31:0]    reg_psum_59_3;
wire signed[31:0]    reg_weight_59_4;
wire signed[31:0]    reg_psum_59_4;
wire signed[31:0]    reg_weight_59_5;
wire signed[31:0]    reg_psum_59_5;
wire signed[31:0]    reg_weight_59_6;
wire signed[31:0]    reg_psum_59_6;
wire signed[31:0]    reg_weight_59_7;
wire signed[31:0]    reg_psum_59_7;
wire signed[31:0]    reg_weight_59_8;
wire signed[31:0]    reg_psum_59_8;
wire signed[31:0]    reg_weight_59_9;
wire signed[31:0]    reg_psum_59_9;
wire signed[31:0]    reg_weight_59_10;
wire signed[31:0]    reg_psum_59_10;
wire signed[31:0]    reg_weight_59_11;
wire signed[31:0]    reg_psum_59_11;
wire signed[31:0]    reg_weight_59_12;
wire signed[31:0]    reg_psum_59_12;
wire signed[31:0]    reg_weight_59_13;
wire signed[31:0]    reg_psum_59_13;
wire signed[31:0]    reg_weight_59_14;
wire signed[31:0]    reg_psum_59_14;
wire signed[31:0]    reg_weight_59_15;
wire signed[31:0]    reg_psum_59_15;
wire signed[31:0]    reg_weight_59_16;
wire signed[31:0]    reg_psum_59_16;
wire signed[31:0]    reg_weight_59_17;
wire signed[31:0]    reg_psum_59_17;
wire signed[31:0]    reg_weight_59_18;
wire signed[31:0]    reg_psum_59_18;
wire signed[31:0]    reg_weight_59_19;
wire signed[31:0]    reg_psum_59_19;
wire signed[31:0]    reg_weight_59_20;
wire signed[31:0]    reg_psum_59_20;
wire signed[31:0]    reg_weight_59_21;
wire signed[31:0]    reg_psum_59_21;
wire signed[31:0]    reg_weight_59_22;
wire signed[31:0]    reg_psum_59_22;
wire signed[31:0]    reg_weight_59_23;
wire signed[31:0]    reg_psum_59_23;
wire signed[31:0]    reg_weight_59_24;
wire signed[31:0]    reg_psum_59_24;
wire signed[31:0]    reg_weight_59_25;
wire signed[31:0]    reg_psum_59_25;
wire signed[31:0]    reg_weight_59_26;
wire signed[31:0]    reg_psum_59_26;
wire signed[31:0]    reg_weight_59_27;
wire signed[31:0]    reg_psum_59_27;
wire signed[31:0]    reg_weight_59_28;
wire signed[31:0]    reg_psum_59_28;
wire signed[31:0]    reg_weight_59_29;
wire signed[31:0]    reg_psum_59_29;
wire signed[31:0]    reg_weight_59_30;
wire signed[31:0]    reg_psum_59_30;
wire signed[31:0]    reg_weight_59_31;
wire signed[31:0]    reg_psum_59_31;
wire signed[31:0]    reg_weight_59_32;
wire signed[31:0]    reg_psum_59_32;
wire signed[31:0]    reg_weight_59_33;
wire signed[31:0]    reg_psum_59_33;
wire signed[31:0]    reg_weight_59_34;
wire signed[31:0]    reg_psum_59_34;
wire signed[31:0]    reg_weight_59_35;
wire signed[31:0]    reg_psum_59_35;
wire signed[31:0]    reg_weight_59_36;
wire signed[31:0]    reg_psum_59_36;
wire signed[31:0]    reg_weight_59_37;
wire signed[31:0]    reg_psum_59_37;
wire signed[31:0]    reg_weight_59_38;
wire signed[31:0]    reg_psum_59_38;
wire signed[31:0]    reg_weight_59_39;
wire signed[31:0]    reg_psum_59_39;
wire signed[31:0]    reg_weight_59_40;
wire signed[31:0]    reg_psum_59_40;
wire signed[31:0]    reg_weight_59_41;
wire signed[31:0]    reg_psum_59_41;
wire signed[31:0]    reg_weight_59_42;
wire signed[31:0]    reg_psum_59_42;
wire signed[31:0]    reg_weight_59_43;
wire signed[31:0]    reg_psum_59_43;
wire signed[31:0]    reg_weight_59_44;
wire signed[31:0]    reg_psum_59_44;
wire signed[31:0]    reg_weight_59_45;
wire signed[31:0]    reg_psum_59_45;
wire signed[31:0]    reg_weight_59_46;
wire signed[31:0]    reg_psum_59_46;
wire signed[31:0]    reg_weight_59_47;
wire signed[31:0]    reg_psum_59_47;
wire signed[31:0]    reg_weight_59_48;
wire signed[31:0]    reg_psum_59_48;
wire signed[31:0]    reg_weight_59_49;
wire signed[31:0]    reg_psum_59_49;
wire signed[31:0]    reg_weight_59_50;
wire signed[31:0]    reg_psum_59_50;
wire signed[31:0]    reg_weight_59_51;
wire signed[31:0]    reg_psum_59_51;
wire signed[31:0]    reg_weight_59_52;
wire signed[31:0]    reg_psum_59_52;
wire signed[31:0]    reg_weight_59_53;
wire signed[31:0]    reg_psum_59_53;
wire signed[31:0]    reg_weight_59_54;
wire signed[31:0]    reg_psum_59_54;
wire signed[31:0]    reg_weight_59_55;
wire signed[31:0]    reg_psum_59_55;
wire signed[31:0]    reg_weight_59_56;
wire signed[31:0]    reg_psum_59_56;
wire signed[31:0]    reg_weight_59_57;
wire signed[31:0]    reg_psum_59_57;
wire signed[31:0]    reg_weight_59_58;
wire signed[31:0]    reg_psum_59_58;
wire signed[31:0]    reg_weight_59_59;
wire signed[31:0]    reg_psum_59_59;
wire signed[31:0]    reg_weight_59_60;
wire signed[31:0]    reg_psum_59_60;
wire signed[31:0]    reg_weight_59_61;
wire signed[31:0]    reg_psum_59_61;
wire signed[31:0]    reg_weight_59_62;
wire signed[31:0]    reg_psum_59_62;
wire signed[31:0]    reg_weight_59_63;
wire signed[31:0]    reg_psum_59_63;
wire signed[31:0]    reg_weight_60_0;
wire signed[31:0]    reg_psum_60_0;
wire signed[31:0]    reg_weight_60_1;
wire signed[31:0]    reg_psum_60_1;
wire signed[31:0]    reg_weight_60_2;
wire signed[31:0]    reg_psum_60_2;
wire signed[31:0]    reg_weight_60_3;
wire signed[31:0]    reg_psum_60_3;
wire signed[31:0]    reg_weight_60_4;
wire signed[31:0]    reg_psum_60_4;
wire signed[31:0]    reg_weight_60_5;
wire signed[31:0]    reg_psum_60_5;
wire signed[31:0]    reg_weight_60_6;
wire signed[31:0]    reg_psum_60_6;
wire signed[31:0]    reg_weight_60_7;
wire signed[31:0]    reg_psum_60_7;
wire signed[31:0]    reg_weight_60_8;
wire signed[31:0]    reg_psum_60_8;
wire signed[31:0]    reg_weight_60_9;
wire signed[31:0]    reg_psum_60_9;
wire signed[31:0]    reg_weight_60_10;
wire signed[31:0]    reg_psum_60_10;
wire signed[31:0]    reg_weight_60_11;
wire signed[31:0]    reg_psum_60_11;
wire signed[31:0]    reg_weight_60_12;
wire signed[31:0]    reg_psum_60_12;
wire signed[31:0]    reg_weight_60_13;
wire signed[31:0]    reg_psum_60_13;
wire signed[31:0]    reg_weight_60_14;
wire signed[31:0]    reg_psum_60_14;
wire signed[31:0]    reg_weight_60_15;
wire signed[31:0]    reg_psum_60_15;
wire signed[31:0]    reg_weight_60_16;
wire signed[31:0]    reg_psum_60_16;
wire signed[31:0]    reg_weight_60_17;
wire signed[31:0]    reg_psum_60_17;
wire signed[31:0]    reg_weight_60_18;
wire signed[31:0]    reg_psum_60_18;
wire signed[31:0]    reg_weight_60_19;
wire signed[31:0]    reg_psum_60_19;
wire signed[31:0]    reg_weight_60_20;
wire signed[31:0]    reg_psum_60_20;
wire signed[31:0]    reg_weight_60_21;
wire signed[31:0]    reg_psum_60_21;
wire signed[31:0]    reg_weight_60_22;
wire signed[31:0]    reg_psum_60_22;
wire signed[31:0]    reg_weight_60_23;
wire signed[31:0]    reg_psum_60_23;
wire signed[31:0]    reg_weight_60_24;
wire signed[31:0]    reg_psum_60_24;
wire signed[31:0]    reg_weight_60_25;
wire signed[31:0]    reg_psum_60_25;
wire signed[31:0]    reg_weight_60_26;
wire signed[31:0]    reg_psum_60_26;
wire signed[31:0]    reg_weight_60_27;
wire signed[31:0]    reg_psum_60_27;
wire signed[31:0]    reg_weight_60_28;
wire signed[31:0]    reg_psum_60_28;
wire signed[31:0]    reg_weight_60_29;
wire signed[31:0]    reg_psum_60_29;
wire signed[31:0]    reg_weight_60_30;
wire signed[31:0]    reg_psum_60_30;
wire signed[31:0]    reg_weight_60_31;
wire signed[31:0]    reg_psum_60_31;
wire signed[31:0]    reg_weight_60_32;
wire signed[31:0]    reg_psum_60_32;
wire signed[31:0]    reg_weight_60_33;
wire signed[31:0]    reg_psum_60_33;
wire signed[31:0]    reg_weight_60_34;
wire signed[31:0]    reg_psum_60_34;
wire signed[31:0]    reg_weight_60_35;
wire signed[31:0]    reg_psum_60_35;
wire signed[31:0]    reg_weight_60_36;
wire signed[31:0]    reg_psum_60_36;
wire signed[31:0]    reg_weight_60_37;
wire signed[31:0]    reg_psum_60_37;
wire signed[31:0]    reg_weight_60_38;
wire signed[31:0]    reg_psum_60_38;
wire signed[31:0]    reg_weight_60_39;
wire signed[31:0]    reg_psum_60_39;
wire signed[31:0]    reg_weight_60_40;
wire signed[31:0]    reg_psum_60_40;
wire signed[31:0]    reg_weight_60_41;
wire signed[31:0]    reg_psum_60_41;
wire signed[31:0]    reg_weight_60_42;
wire signed[31:0]    reg_psum_60_42;
wire signed[31:0]    reg_weight_60_43;
wire signed[31:0]    reg_psum_60_43;
wire signed[31:0]    reg_weight_60_44;
wire signed[31:0]    reg_psum_60_44;
wire signed[31:0]    reg_weight_60_45;
wire signed[31:0]    reg_psum_60_45;
wire signed[31:0]    reg_weight_60_46;
wire signed[31:0]    reg_psum_60_46;
wire signed[31:0]    reg_weight_60_47;
wire signed[31:0]    reg_psum_60_47;
wire signed[31:0]    reg_weight_60_48;
wire signed[31:0]    reg_psum_60_48;
wire signed[31:0]    reg_weight_60_49;
wire signed[31:0]    reg_psum_60_49;
wire signed[31:0]    reg_weight_60_50;
wire signed[31:0]    reg_psum_60_50;
wire signed[31:0]    reg_weight_60_51;
wire signed[31:0]    reg_psum_60_51;
wire signed[31:0]    reg_weight_60_52;
wire signed[31:0]    reg_psum_60_52;
wire signed[31:0]    reg_weight_60_53;
wire signed[31:0]    reg_psum_60_53;
wire signed[31:0]    reg_weight_60_54;
wire signed[31:0]    reg_psum_60_54;
wire signed[31:0]    reg_weight_60_55;
wire signed[31:0]    reg_psum_60_55;
wire signed[31:0]    reg_weight_60_56;
wire signed[31:0]    reg_psum_60_56;
wire signed[31:0]    reg_weight_60_57;
wire signed[31:0]    reg_psum_60_57;
wire signed[31:0]    reg_weight_60_58;
wire signed[31:0]    reg_psum_60_58;
wire signed[31:0]    reg_weight_60_59;
wire signed[31:0]    reg_psum_60_59;
wire signed[31:0]    reg_weight_60_60;
wire signed[31:0]    reg_psum_60_60;
wire signed[31:0]    reg_weight_60_61;
wire signed[31:0]    reg_psum_60_61;
wire signed[31:0]    reg_weight_60_62;
wire signed[31:0]    reg_psum_60_62;
wire signed[31:0]    reg_weight_60_63;
wire signed[31:0]    reg_psum_60_63;
wire signed[31:0]    reg_weight_61_0;
wire signed[31:0]    reg_psum_61_0;
wire signed[31:0]    reg_weight_61_1;
wire signed[31:0]    reg_psum_61_1;
wire signed[31:0]    reg_weight_61_2;
wire signed[31:0]    reg_psum_61_2;
wire signed[31:0]    reg_weight_61_3;
wire signed[31:0]    reg_psum_61_3;
wire signed[31:0]    reg_weight_61_4;
wire signed[31:0]    reg_psum_61_4;
wire signed[31:0]    reg_weight_61_5;
wire signed[31:0]    reg_psum_61_5;
wire signed[31:0]    reg_weight_61_6;
wire signed[31:0]    reg_psum_61_6;
wire signed[31:0]    reg_weight_61_7;
wire signed[31:0]    reg_psum_61_7;
wire signed[31:0]    reg_weight_61_8;
wire signed[31:0]    reg_psum_61_8;
wire signed[31:0]    reg_weight_61_9;
wire signed[31:0]    reg_psum_61_9;
wire signed[31:0]    reg_weight_61_10;
wire signed[31:0]    reg_psum_61_10;
wire signed[31:0]    reg_weight_61_11;
wire signed[31:0]    reg_psum_61_11;
wire signed[31:0]    reg_weight_61_12;
wire signed[31:0]    reg_psum_61_12;
wire signed[31:0]    reg_weight_61_13;
wire signed[31:0]    reg_psum_61_13;
wire signed[31:0]    reg_weight_61_14;
wire signed[31:0]    reg_psum_61_14;
wire signed[31:0]    reg_weight_61_15;
wire signed[31:0]    reg_psum_61_15;
wire signed[31:0]    reg_weight_61_16;
wire signed[31:0]    reg_psum_61_16;
wire signed[31:0]    reg_weight_61_17;
wire signed[31:0]    reg_psum_61_17;
wire signed[31:0]    reg_weight_61_18;
wire signed[31:0]    reg_psum_61_18;
wire signed[31:0]    reg_weight_61_19;
wire signed[31:0]    reg_psum_61_19;
wire signed[31:0]    reg_weight_61_20;
wire signed[31:0]    reg_psum_61_20;
wire signed[31:0]    reg_weight_61_21;
wire signed[31:0]    reg_psum_61_21;
wire signed[31:0]    reg_weight_61_22;
wire signed[31:0]    reg_psum_61_22;
wire signed[31:0]    reg_weight_61_23;
wire signed[31:0]    reg_psum_61_23;
wire signed[31:0]    reg_weight_61_24;
wire signed[31:0]    reg_psum_61_24;
wire signed[31:0]    reg_weight_61_25;
wire signed[31:0]    reg_psum_61_25;
wire signed[31:0]    reg_weight_61_26;
wire signed[31:0]    reg_psum_61_26;
wire signed[31:0]    reg_weight_61_27;
wire signed[31:0]    reg_psum_61_27;
wire signed[31:0]    reg_weight_61_28;
wire signed[31:0]    reg_psum_61_28;
wire signed[31:0]    reg_weight_61_29;
wire signed[31:0]    reg_psum_61_29;
wire signed[31:0]    reg_weight_61_30;
wire signed[31:0]    reg_psum_61_30;
wire signed[31:0]    reg_weight_61_31;
wire signed[31:0]    reg_psum_61_31;
wire signed[31:0]    reg_weight_61_32;
wire signed[31:0]    reg_psum_61_32;
wire signed[31:0]    reg_weight_61_33;
wire signed[31:0]    reg_psum_61_33;
wire signed[31:0]    reg_weight_61_34;
wire signed[31:0]    reg_psum_61_34;
wire signed[31:0]    reg_weight_61_35;
wire signed[31:0]    reg_psum_61_35;
wire signed[31:0]    reg_weight_61_36;
wire signed[31:0]    reg_psum_61_36;
wire signed[31:0]    reg_weight_61_37;
wire signed[31:0]    reg_psum_61_37;
wire signed[31:0]    reg_weight_61_38;
wire signed[31:0]    reg_psum_61_38;
wire signed[31:0]    reg_weight_61_39;
wire signed[31:0]    reg_psum_61_39;
wire signed[31:0]    reg_weight_61_40;
wire signed[31:0]    reg_psum_61_40;
wire signed[31:0]    reg_weight_61_41;
wire signed[31:0]    reg_psum_61_41;
wire signed[31:0]    reg_weight_61_42;
wire signed[31:0]    reg_psum_61_42;
wire signed[31:0]    reg_weight_61_43;
wire signed[31:0]    reg_psum_61_43;
wire signed[31:0]    reg_weight_61_44;
wire signed[31:0]    reg_psum_61_44;
wire signed[31:0]    reg_weight_61_45;
wire signed[31:0]    reg_psum_61_45;
wire signed[31:0]    reg_weight_61_46;
wire signed[31:0]    reg_psum_61_46;
wire signed[31:0]    reg_weight_61_47;
wire signed[31:0]    reg_psum_61_47;
wire signed[31:0]    reg_weight_61_48;
wire signed[31:0]    reg_psum_61_48;
wire signed[31:0]    reg_weight_61_49;
wire signed[31:0]    reg_psum_61_49;
wire signed[31:0]    reg_weight_61_50;
wire signed[31:0]    reg_psum_61_50;
wire signed[31:0]    reg_weight_61_51;
wire signed[31:0]    reg_psum_61_51;
wire signed[31:0]    reg_weight_61_52;
wire signed[31:0]    reg_psum_61_52;
wire signed[31:0]    reg_weight_61_53;
wire signed[31:0]    reg_psum_61_53;
wire signed[31:0]    reg_weight_61_54;
wire signed[31:0]    reg_psum_61_54;
wire signed[31:0]    reg_weight_61_55;
wire signed[31:0]    reg_psum_61_55;
wire signed[31:0]    reg_weight_61_56;
wire signed[31:0]    reg_psum_61_56;
wire signed[31:0]    reg_weight_61_57;
wire signed[31:0]    reg_psum_61_57;
wire signed[31:0]    reg_weight_61_58;
wire signed[31:0]    reg_psum_61_58;
wire signed[31:0]    reg_weight_61_59;
wire signed[31:0]    reg_psum_61_59;
wire signed[31:0]    reg_weight_61_60;
wire signed[31:0]    reg_psum_61_60;
wire signed[31:0]    reg_weight_61_61;
wire signed[31:0]    reg_psum_61_61;
wire signed[31:0]    reg_weight_61_62;
wire signed[31:0]    reg_psum_61_62;
wire signed[31:0]    reg_weight_61_63;
wire signed[31:0]    reg_psum_61_63;
wire signed[31:0]    reg_weight_62_0;
wire signed[31:0]    reg_psum_62_0;
wire signed[31:0]    reg_weight_62_1;
wire signed[31:0]    reg_psum_62_1;
wire signed[31:0]    reg_weight_62_2;
wire signed[31:0]    reg_psum_62_2;
wire signed[31:0]    reg_weight_62_3;
wire signed[31:0]    reg_psum_62_3;
wire signed[31:0]    reg_weight_62_4;
wire signed[31:0]    reg_psum_62_4;
wire signed[31:0]    reg_weight_62_5;
wire signed[31:0]    reg_psum_62_5;
wire signed[31:0]    reg_weight_62_6;
wire signed[31:0]    reg_psum_62_6;
wire signed[31:0]    reg_weight_62_7;
wire signed[31:0]    reg_psum_62_7;
wire signed[31:0]    reg_weight_62_8;
wire signed[31:0]    reg_psum_62_8;
wire signed[31:0]    reg_weight_62_9;
wire signed[31:0]    reg_psum_62_9;
wire signed[31:0]    reg_weight_62_10;
wire signed[31:0]    reg_psum_62_10;
wire signed[31:0]    reg_weight_62_11;
wire signed[31:0]    reg_psum_62_11;
wire signed[31:0]    reg_weight_62_12;
wire signed[31:0]    reg_psum_62_12;
wire signed[31:0]    reg_weight_62_13;
wire signed[31:0]    reg_psum_62_13;
wire signed[31:0]    reg_weight_62_14;
wire signed[31:0]    reg_psum_62_14;
wire signed[31:0]    reg_weight_62_15;
wire signed[31:0]    reg_psum_62_15;
wire signed[31:0]    reg_weight_62_16;
wire signed[31:0]    reg_psum_62_16;
wire signed[31:0]    reg_weight_62_17;
wire signed[31:0]    reg_psum_62_17;
wire signed[31:0]    reg_weight_62_18;
wire signed[31:0]    reg_psum_62_18;
wire signed[31:0]    reg_weight_62_19;
wire signed[31:0]    reg_psum_62_19;
wire signed[31:0]    reg_weight_62_20;
wire signed[31:0]    reg_psum_62_20;
wire signed[31:0]    reg_weight_62_21;
wire signed[31:0]    reg_psum_62_21;
wire signed[31:0]    reg_weight_62_22;
wire signed[31:0]    reg_psum_62_22;
wire signed[31:0]    reg_weight_62_23;
wire signed[31:0]    reg_psum_62_23;
wire signed[31:0]    reg_weight_62_24;
wire signed[31:0]    reg_psum_62_24;
wire signed[31:0]    reg_weight_62_25;
wire signed[31:0]    reg_psum_62_25;
wire signed[31:0]    reg_weight_62_26;
wire signed[31:0]    reg_psum_62_26;
wire signed[31:0]    reg_weight_62_27;
wire signed[31:0]    reg_psum_62_27;
wire signed[31:0]    reg_weight_62_28;
wire signed[31:0]    reg_psum_62_28;
wire signed[31:0]    reg_weight_62_29;
wire signed[31:0]    reg_psum_62_29;
wire signed[31:0]    reg_weight_62_30;
wire signed[31:0]    reg_psum_62_30;
wire signed[31:0]    reg_weight_62_31;
wire signed[31:0]    reg_psum_62_31;
wire signed[31:0]    reg_weight_62_32;
wire signed[31:0]    reg_psum_62_32;
wire signed[31:0]    reg_weight_62_33;
wire signed[31:0]    reg_psum_62_33;
wire signed[31:0]    reg_weight_62_34;
wire signed[31:0]    reg_psum_62_34;
wire signed[31:0]    reg_weight_62_35;
wire signed[31:0]    reg_psum_62_35;
wire signed[31:0]    reg_weight_62_36;
wire signed[31:0]    reg_psum_62_36;
wire signed[31:0]    reg_weight_62_37;
wire signed[31:0]    reg_psum_62_37;
wire signed[31:0]    reg_weight_62_38;
wire signed[31:0]    reg_psum_62_38;
wire signed[31:0]    reg_weight_62_39;
wire signed[31:0]    reg_psum_62_39;
wire signed[31:0]    reg_weight_62_40;
wire signed[31:0]    reg_psum_62_40;
wire signed[31:0]    reg_weight_62_41;
wire signed[31:0]    reg_psum_62_41;
wire signed[31:0]    reg_weight_62_42;
wire signed[31:0]    reg_psum_62_42;
wire signed[31:0]    reg_weight_62_43;
wire signed[31:0]    reg_psum_62_43;
wire signed[31:0]    reg_weight_62_44;
wire signed[31:0]    reg_psum_62_44;
wire signed[31:0]    reg_weight_62_45;
wire signed[31:0]    reg_psum_62_45;
wire signed[31:0]    reg_weight_62_46;
wire signed[31:0]    reg_psum_62_46;
wire signed[31:0]    reg_weight_62_47;
wire signed[31:0]    reg_psum_62_47;
wire signed[31:0]    reg_weight_62_48;
wire signed[31:0]    reg_psum_62_48;
wire signed[31:0]    reg_weight_62_49;
wire signed[31:0]    reg_psum_62_49;
wire signed[31:0]    reg_weight_62_50;
wire signed[31:0]    reg_psum_62_50;
wire signed[31:0]    reg_weight_62_51;
wire signed[31:0]    reg_psum_62_51;
wire signed[31:0]    reg_weight_62_52;
wire signed[31:0]    reg_psum_62_52;
wire signed[31:0]    reg_weight_62_53;
wire signed[31:0]    reg_psum_62_53;
wire signed[31:0]    reg_weight_62_54;
wire signed[31:0]    reg_psum_62_54;
wire signed[31:0]    reg_weight_62_55;
wire signed[31:0]    reg_psum_62_55;
wire signed[31:0]    reg_weight_62_56;
wire signed[31:0]    reg_psum_62_56;
wire signed[31:0]    reg_weight_62_57;
wire signed[31:0]    reg_psum_62_57;
wire signed[31:0]    reg_weight_62_58;
wire signed[31:0]    reg_psum_62_58;
wire signed[31:0]    reg_weight_62_59;
wire signed[31:0]    reg_psum_62_59;
wire signed[31:0]    reg_weight_62_60;
wire signed[31:0]    reg_psum_62_60;
wire signed[31:0]    reg_weight_62_61;
wire signed[31:0]    reg_psum_62_61;
wire signed[31:0]    reg_weight_62_62;
wire signed[31:0]    reg_psum_62_62;
wire signed[31:0]    reg_weight_62_63;
wire signed[31:0]    reg_psum_62_63;
wire signed[31:0]    reg_weight_63_0;
wire signed[31:0]    reg_psum_63_0;
wire signed[31:0]    reg_weight_63_1;
wire signed[31:0]    reg_psum_63_1;
wire signed[31:0]    reg_weight_63_2;
wire signed[31:0]    reg_psum_63_2;
wire signed[31:0]    reg_weight_63_3;
wire signed[31:0]    reg_psum_63_3;
wire signed[31:0]    reg_weight_63_4;
wire signed[31:0]    reg_psum_63_4;
wire signed[31:0]    reg_weight_63_5;
wire signed[31:0]    reg_psum_63_5;
wire signed[31:0]    reg_weight_63_6;
wire signed[31:0]    reg_psum_63_6;
wire signed[31:0]    reg_weight_63_7;
wire signed[31:0]    reg_psum_63_7;
wire signed[31:0]    reg_weight_63_8;
wire signed[31:0]    reg_psum_63_8;
wire signed[31:0]    reg_weight_63_9;
wire signed[31:0]    reg_psum_63_9;
wire signed[31:0]    reg_weight_63_10;
wire signed[31:0]    reg_psum_63_10;
wire signed[31:0]    reg_weight_63_11;
wire signed[31:0]    reg_psum_63_11;
wire signed[31:0]    reg_weight_63_12;
wire signed[31:0]    reg_psum_63_12;
wire signed[31:0]    reg_weight_63_13;
wire signed[31:0]    reg_psum_63_13;
wire signed[31:0]    reg_weight_63_14;
wire signed[31:0]    reg_psum_63_14;
wire signed[31:0]    reg_weight_63_15;
wire signed[31:0]    reg_psum_63_15;
wire signed[31:0]    reg_weight_63_16;
wire signed[31:0]    reg_psum_63_16;
wire signed[31:0]    reg_weight_63_17;
wire signed[31:0]    reg_psum_63_17;
wire signed[31:0]    reg_weight_63_18;
wire signed[31:0]    reg_psum_63_18;
wire signed[31:0]    reg_weight_63_19;
wire signed[31:0]    reg_psum_63_19;
wire signed[31:0]    reg_weight_63_20;
wire signed[31:0]    reg_psum_63_20;
wire signed[31:0]    reg_weight_63_21;
wire signed[31:0]    reg_psum_63_21;
wire signed[31:0]    reg_weight_63_22;
wire signed[31:0]    reg_psum_63_22;
wire signed[31:0]    reg_weight_63_23;
wire signed[31:0]    reg_psum_63_23;
wire signed[31:0]    reg_weight_63_24;
wire signed[31:0]    reg_psum_63_24;
wire signed[31:0]    reg_weight_63_25;
wire signed[31:0]    reg_psum_63_25;
wire signed[31:0]    reg_weight_63_26;
wire signed[31:0]    reg_psum_63_26;
wire signed[31:0]    reg_weight_63_27;
wire signed[31:0]    reg_psum_63_27;
wire signed[31:0]    reg_weight_63_28;
wire signed[31:0]    reg_psum_63_28;
wire signed[31:0]    reg_weight_63_29;
wire signed[31:0]    reg_psum_63_29;
wire signed[31:0]    reg_weight_63_30;
wire signed[31:0]    reg_psum_63_30;
wire signed[31:0]    reg_weight_63_31;
wire signed[31:0]    reg_psum_63_31;
wire signed[31:0]    reg_weight_63_32;
wire signed[31:0]    reg_psum_63_32;
wire signed[31:0]    reg_weight_63_33;
wire signed[31:0]    reg_psum_63_33;
wire signed[31:0]    reg_weight_63_34;
wire signed[31:0]    reg_psum_63_34;
wire signed[31:0]    reg_weight_63_35;
wire signed[31:0]    reg_psum_63_35;
wire signed[31:0]    reg_weight_63_36;
wire signed[31:0]    reg_psum_63_36;
wire signed[31:0]    reg_weight_63_37;
wire signed[31:0]    reg_psum_63_37;
wire signed[31:0]    reg_weight_63_38;
wire signed[31:0]    reg_psum_63_38;
wire signed[31:0]    reg_weight_63_39;
wire signed[31:0]    reg_psum_63_39;
wire signed[31:0]    reg_weight_63_40;
wire signed[31:0]    reg_psum_63_40;
wire signed[31:0]    reg_weight_63_41;
wire signed[31:0]    reg_psum_63_41;
wire signed[31:0]    reg_weight_63_42;
wire signed[31:0]    reg_psum_63_42;
wire signed[31:0]    reg_weight_63_43;
wire signed[31:0]    reg_psum_63_43;
wire signed[31:0]    reg_weight_63_44;
wire signed[31:0]    reg_psum_63_44;
wire signed[31:0]    reg_weight_63_45;
wire signed[31:0]    reg_psum_63_45;
wire signed[31:0]    reg_weight_63_46;
wire signed[31:0]    reg_psum_63_46;
wire signed[31:0]    reg_weight_63_47;
wire signed[31:0]    reg_psum_63_47;
wire signed[31:0]    reg_weight_63_48;
wire signed[31:0]    reg_psum_63_48;
wire signed[31:0]    reg_weight_63_49;
wire signed[31:0]    reg_psum_63_49;
wire signed[31:0]    reg_weight_63_50;
wire signed[31:0]    reg_psum_63_50;
wire signed[31:0]    reg_weight_63_51;
wire signed[31:0]    reg_psum_63_51;
wire signed[31:0]    reg_weight_63_52;
wire signed[31:0]    reg_psum_63_52;
wire signed[31:0]    reg_weight_63_53;
wire signed[31:0]    reg_psum_63_53;
wire signed[31:0]    reg_weight_63_54;
wire signed[31:0]    reg_psum_63_54;
wire signed[31:0]    reg_weight_63_55;
wire signed[31:0]    reg_psum_63_55;
wire signed[31:0]    reg_weight_63_56;
wire signed[31:0]    reg_psum_63_56;
wire signed[31:0]    reg_weight_63_57;
wire signed[31:0]    reg_psum_63_57;
wire signed[31:0]    reg_weight_63_58;
wire signed[31:0]    reg_psum_63_58;
wire signed[31:0]    reg_weight_63_59;
wire signed[31:0]    reg_psum_63_59;
wire signed[31:0]    reg_weight_63_60;
wire signed[31:0]    reg_psum_63_60;
wire signed[31:0]    reg_weight_63_61;
wire signed[31:0]    reg_psum_63_61;
wire signed[31:0]    reg_weight_63_62;
wire signed[31:0]    reg_psum_63_62;
wire signed[31:0]    reg_weight_63_63;
wire signed[31:0]    reg_psum_63_63;
PE U0_0( .activation_in(in_activation_0), .weight_in(in_weight_0), .partial_sum_in(in_psum_0), .reg_activation(reg_activation_0_0), .reg_weight(reg_weight_0_0), .reg_partial_sum(reg_psum_0_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_1( .activation_in(reg_activation_0_0), .weight_in(in_weight_1), .partial_sum_in(in_psum_1), .reg_activation(reg_activation_0_1), .reg_weight(reg_weight_0_1), .reg_partial_sum(reg_psum_0_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_2( .activation_in(reg_activation_0_1), .weight_in(in_weight_2), .partial_sum_in(in_psum_2), .reg_activation(reg_activation_0_2), .reg_weight(reg_weight_0_2), .reg_partial_sum(reg_psum_0_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_3( .activation_in(reg_activation_0_2), .weight_in(in_weight_3), .partial_sum_in(in_psum_3), .reg_activation(reg_activation_0_3), .reg_weight(reg_weight_0_3), .reg_partial_sum(reg_psum_0_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_4( .activation_in(reg_activation_0_3), .weight_in(in_weight_4), .partial_sum_in(in_psum_4), .reg_activation(reg_activation_0_4), .reg_weight(reg_weight_0_4), .reg_partial_sum(reg_psum_0_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_5( .activation_in(reg_activation_0_4), .weight_in(in_weight_5), .partial_sum_in(in_psum_5), .reg_activation(reg_activation_0_5), .reg_weight(reg_weight_0_5), .reg_partial_sum(reg_psum_0_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_6( .activation_in(reg_activation_0_5), .weight_in(in_weight_6), .partial_sum_in(in_psum_6), .reg_activation(reg_activation_0_6), .reg_weight(reg_weight_0_6), .reg_partial_sum(reg_psum_0_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_7( .activation_in(reg_activation_0_6), .weight_in(in_weight_7), .partial_sum_in(in_psum_7), .reg_activation(reg_activation_0_7), .reg_weight(reg_weight_0_7), .reg_partial_sum(reg_psum_0_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_8( .activation_in(reg_activation_0_7), .weight_in(in_weight_8), .partial_sum_in(in_psum_8), .reg_activation(reg_activation_0_8), .reg_weight(reg_weight_0_8), .reg_partial_sum(reg_psum_0_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_9( .activation_in(reg_activation_0_8), .weight_in(in_weight_9), .partial_sum_in(in_psum_9), .reg_activation(reg_activation_0_9), .reg_weight(reg_weight_0_9), .reg_partial_sum(reg_psum_0_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_10( .activation_in(reg_activation_0_9), .weight_in(in_weight_10), .partial_sum_in(in_psum_10), .reg_activation(reg_activation_0_10), .reg_weight(reg_weight_0_10), .reg_partial_sum(reg_psum_0_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_11( .activation_in(reg_activation_0_10), .weight_in(in_weight_11), .partial_sum_in(in_psum_11), .reg_activation(reg_activation_0_11), .reg_weight(reg_weight_0_11), .reg_partial_sum(reg_psum_0_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_12( .activation_in(reg_activation_0_11), .weight_in(in_weight_12), .partial_sum_in(in_psum_12), .reg_activation(reg_activation_0_12), .reg_weight(reg_weight_0_12), .reg_partial_sum(reg_psum_0_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_13( .activation_in(reg_activation_0_12), .weight_in(in_weight_13), .partial_sum_in(in_psum_13), .reg_activation(reg_activation_0_13), .reg_weight(reg_weight_0_13), .reg_partial_sum(reg_psum_0_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_14( .activation_in(reg_activation_0_13), .weight_in(in_weight_14), .partial_sum_in(in_psum_14), .reg_activation(reg_activation_0_14), .reg_weight(reg_weight_0_14), .reg_partial_sum(reg_psum_0_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_15( .activation_in(reg_activation_0_14), .weight_in(in_weight_15), .partial_sum_in(in_psum_15), .reg_activation(reg_activation_0_15), .reg_weight(reg_weight_0_15), .reg_partial_sum(reg_psum_0_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_16( .activation_in(reg_activation_0_15), .weight_in(in_weight_16), .partial_sum_in(in_psum_16), .reg_activation(reg_activation_0_16), .reg_weight(reg_weight_0_16), .reg_partial_sum(reg_psum_0_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_17( .activation_in(reg_activation_0_16), .weight_in(in_weight_17), .partial_sum_in(in_psum_17), .reg_activation(reg_activation_0_17), .reg_weight(reg_weight_0_17), .reg_partial_sum(reg_psum_0_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_18( .activation_in(reg_activation_0_17), .weight_in(in_weight_18), .partial_sum_in(in_psum_18), .reg_activation(reg_activation_0_18), .reg_weight(reg_weight_0_18), .reg_partial_sum(reg_psum_0_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_19( .activation_in(reg_activation_0_18), .weight_in(in_weight_19), .partial_sum_in(in_psum_19), .reg_activation(reg_activation_0_19), .reg_weight(reg_weight_0_19), .reg_partial_sum(reg_psum_0_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_20( .activation_in(reg_activation_0_19), .weight_in(in_weight_20), .partial_sum_in(in_psum_20), .reg_activation(reg_activation_0_20), .reg_weight(reg_weight_0_20), .reg_partial_sum(reg_psum_0_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_21( .activation_in(reg_activation_0_20), .weight_in(in_weight_21), .partial_sum_in(in_psum_21), .reg_activation(reg_activation_0_21), .reg_weight(reg_weight_0_21), .reg_partial_sum(reg_psum_0_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_22( .activation_in(reg_activation_0_21), .weight_in(in_weight_22), .partial_sum_in(in_psum_22), .reg_activation(reg_activation_0_22), .reg_weight(reg_weight_0_22), .reg_partial_sum(reg_psum_0_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_23( .activation_in(reg_activation_0_22), .weight_in(in_weight_23), .partial_sum_in(in_psum_23), .reg_activation(reg_activation_0_23), .reg_weight(reg_weight_0_23), .reg_partial_sum(reg_psum_0_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_24( .activation_in(reg_activation_0_23), .weight_in(in_weight_24), .partial_sum_in(in_psum_24), .reg_activation(reg_activation_0_24), .reg_weight(reg_weight_0_24), .reg_partial_sum(reg_psum_0_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_25( .activation_in(reg_activation_0_24), .weight_in(in_weight_25), .partial_sum_in(in_psum_25), .reg_activation(reg_activation_0_25), .reg_weight(reg_weight_0_25), .reg_partial_sum(reg_psum_0_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_26( .activation_in(reg_activation_0_25), .weight_in(in_weight_26), .partial_sum_in(in_psum_26), .reg_activation(reg_activation_0_26), .reg_weight(reg_weight_0_26), .reg_partial_sum(reg_psum_0_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_27( .activation_in(reg_activation_0_26), .weight_in(in_weight_27), .partial_sum_in(in_psum_27), .reg_activation(reg_activation_0_27), .reg_weight(reg_weight_0_27), .reg_partial_sum(reg_psum_0_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_28( .activation_in(reg_activation_0_27), .weight_in(in_weight_28), .partial_sum_in(in_psum_28), .reg_activation(reg_activation_0_28), .reg_weight(reg_weight_0_28), .reg_partial_sum(reg_psum_0_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_29( .activation_in(reg_activation_0_28), .weight_in(in_weight_29), .partial_sum_in(in_psum_29), .reg_activation(reg_activation_0_29), .reg_weight(reg_weight_0_29), .reg_partial_sum(reg_psum_0_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_30( .activation_in(reg_activation_0_29), .weight_in(in_weight_30), .partial_sum_in(in_psum_30), .reg_activation(reg_activation_0_30), .reg_weight(reg_weight_0_30), .reg_partial_sum(reg_psum_0_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_31( .activation_in(reg_activation_0_30), .weight_in(in_weight_31), .partial_sum_in(in_psum_31), .reg_activation(reg_activation_0_31), .reg_weight(reg_weight_0_31), .reg_partial_sum(reg_psum_0_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_32( .activation_in(reg_activation_0_31), .weight_in(in_weight_32), .partial_sum_in(in_psum_32), .reg_activation(reg_activation_0_32), .reg_weight(reg_weight_0_32), .reg_partial_sum(reg_psum_0_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_33( .activation_in(reg_activation_0_32), .weight_in(in_weight_33), .partial_sum_in(in_psum_33), .reg_activation(reg_activation_0_33), .reg_weight(reg_weight_0_33), .reg_partial_sum(reg_psum_0_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_34( .activation_in(reg_activation_0_33), .weight_in(in_weight_34), .partial_sum_in(in_psum_34), .reg_activation(reg_activation_0_34), .reg_weight(reg_weight_0_34), .reg_partial_sum(reg_psum_0_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_35( .activation_in(reg_activation_0_34), .weight_in(in_weight_35), .partial_sum_in(in_psum_35), .reg_activation(reg_activation_0_35), .reg_weight(reg_weight_0_35), .reg_partial_sum(reg_psum_0_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_36( .activation_in(reg_activation_0_35), .weight_in(in_weight_36), .partial_sum_in(in_psum_36), .reg_activation(reg_activation_0_36), .reg_weight(reg_weight_0_36), .reg_partial_sum(reg_psum_0_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_37( .activation_in(reg_activation_0_36), .weight_in(in_weight_37), .partial_sum_in(in_psum_37), .reg_activation(reg_activation_0_37), .reg_weight(reg_weight_0_37), .reg_partial_sum(reg_psum_0_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_38( .activation_in(reg_activation_0_37), .weight_in(in_weight_38), .partial_sum_in(in_psum_38), .reg_activation(reg_activation_0_38), .reg_weight(reg_weight_0_38), .reg_partial_sum(reg_psum_0_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_39( .activation_in(reg_activation_0_38), .weight_in(in_weight_39), .partial_sum_in(in_psum_39), .reg_activation(reg_activation_0_39), .reg_weight(reg_weight_0_39), .reg_partial_sum(reg_psum_0_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_40( .activation_in(reg_activation_0_39), .weight_in(in_weight_40), .partial_sum_in(in_psum_40), .reg_activation(reg_activation_0_40), .reg_weight(reg_weight_0_40), .reg_partial_sum(reg_psum_0_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_41( .activation_in(reg_activation_0_40), .weight_in(in_weight_41), .partial_sum_in(in_psum_41), .reg_activation(reg_activation_0_41), .reg_weight(reg_weight_0_41), .reg_partial_sum(reg_psum_0_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_42( .activation_in(reg_activation_0_41), .weight_in(in_weight_42), .partial_sum_in(in_psum_42), .reg_activation(reg_activation_0_42), .reg_weight(reg_weight_0_42), .reg_partial_sum(reg_psum_0_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_43( .activation_in(reg_activation_0_42), .weight_in(in_weight_43), .partial_sum_in(in_psum_43), .reg_activation(reg_activation_0_43), .reg_weight(reg_weight_0_43), .reg_partial_sum(reg_psum_0_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_44( .activation_in(reg_activation_0_43), .weight_in(in_weight_44), .partial_sum_in(in_psum_44), .reg_activation(reg_activation_0_44), .reg_weight(reg_weight_0_44), .reg_partial_sum(reg_psum_0_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_45( .activation_in(reg_activation_0_44), .weight_in(in_weight_45), .partial_sum_in(in_psum_45), .reg_activation(reg_activation_0_45), .reg_weight(reg_weight_0_45), .reg_partial_sum(reg_psum_0_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_46( .activation_in(reg_activation_0_45), .weight_in(in_weight_46), .partial_sum_in(in_psum_46), .reg_activation(reg_activation_0_46), .reg_weight(reg_weight_0_46), .reg_partial_sum(reg_psum_0_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_47( .activation_in(reg_activation_0_46), .weight_in(in_weight_47), .partial_sum_in(in_psum_47), .reg_activation(reg_activation_0_47), .reg_weight(reg_weight_0_47), .reg_partial_sum(reg_psum_0_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_48( .activation_in(reg_activation_0_47), .weight_in(in_weight_48), .partial_sum_in(in_psum_48), .reg_activation(reg_activation_0_48), .reg_weight(reg_weight_0_48), .reg_partial_sum(reg_psum_0_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_49( .activation_in(reg_activation_0_48), .weight_in(in_weight_49), .partial_sum_in(in_psum_49), .reg_activation(reg_activation_0_49), .reg_weight(reg_weight_0_49), .reg_partial_sum(reg_psum_0_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_50( .activation_in(reg_activation_0_49), .weight_in(in_weight_50), .partial_sum_in(in_psum_50), .reg_activation(reg_activation_0_50), .reg_weight(reg_weight_0_50), .reg_partial_sum(reg_psum_0_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_51( .activation_in(reg_activation_0_50), .weight_in(in_weight_51), .partial_sum_in(in_psum_51), .reg_activation(reg_activation_0_51), .reg_weight(reg_weight_0_51), .reg_partial_sum(reg_psum_0_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_52( .activation_in(reg_activation_0_51), .weight_in(in_weight_52), .partial_sum_in(in_psum_52), .reg_activation(reg_activation_0_52), .reg_weight(reg_weight_0_52), .reg_partial_sum(reg_psum_0_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_53( .activation_in(reg_activation_0_52), .weight_in(in_weight_53), .partial_sum_in(in_psum_53), .reg_activation(reg_activation_0_53), .reg_weight(reg_weight_0_53), .reg_partial_sum(reg_psum_0_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_54( .activation_in(reg_activation_0_53), .weight_in(in_weight_54), .partial_sum_in(in_psum_54), .reg_activation(reg_activation_0_54), .reg_weight(reg_weight_0_54), .reg_partial_sum(reg_psum_0_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_55( .activation_in(reg_activation_0_54), .weight_in(in_weight_55), .partial_sum_in(in_psum_55), .reg_activation(reg_activation_0_55), .reg_weight(reg_weight_0_55), .reg_partial_sum(reg_psum_0_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_56( .activation_in(reg_activation_0_55), .weight_in(in_weight_56), .partial_sum_in(in_psum_56), .reg_activation(reg_activation_0_56), .reg_weight(reg_weight_0_56), .reg_partial_sum(reg_psum_0_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_57( .activation_in(reg_activation_0_56), .weight_in(in_weight_57), .partial_sum_in(in_psum_57), .reg_activation(reg_activation_0_57), .reg_weight(reg_weight_0_57), .reg_partial_sum(reg_psum_0_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_58( .activation_in(reg_activation_0_57), .weight_in(in_weight_58), .partial_sum_in(in_psum_58), .reg_activation(reg_activation_0_58), .reg_weight(reg_weight_0_58), .reg_partial_sum(reg_psum_0_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_59( .activation_in(reg_activation_0_58), .weight_in(in_weight_59), .partial_sum_in(in_psum_59), .reg_activation(reg_activation_0_59), .reg_weight(reg_weight_0_59), .reg_partial_sum(reg_psum_0_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_60( .activation_in(reg_activation_0_59), .weight_in(in_weight_60), .partial_sum_in(in_psum_60), .reg_activation(reg_activation_0_60), .reg_weight(reg_weight_0_60), .reg_partial_sum(reg_psum_0_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_61( .activation_in(reg_activation_0_60), .weight_in(in_weight_61), .partial_sum_in(in_psum_61), .reg_activation(reg_activation_0_61), .reg_weight(reg_weight_0_61), .reg_partial_sum(reg_psum_0_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_62( .activation_in(reg_activation_0_61), .weight_in(in_weight_62), .partial_sum_in(in_psum_62), .reg_activation(reg_activation_0_62), .reg_weight(reg_weight_0_62), .reg_partial_sum(reg_psum_0_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_63( .activation_in(reg_activation_0_62), .weight_in(in_weight_63), .partial_sum_in(in_psum_63), .reg_weight(reg_weight_0_63), .reg_partial_sum(reg_psum_0_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_0( .activation_in(in_activation_1), .weight_in(reg_weight_0_0), .partial_sum_in(reg_psum_0_0), .reg_activation(reg_activation_1_0), .reg_weight(reg_weight_1_0), .reg_partial_sum(reg_psum_1_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_1( .activation_in(reg_activation_1_0), .weight_in(reg_weight_0_1), .partial_sum_in(reg_psum_0_1), .reg_activation(reg_activation_1_1), .reg_weight(reg_weight_1_1), .reg_partial_sum(reg_psum_1_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_2( .activation_in(reg_activation_1_1), .weight_in(reg_weight_0_2), .partial_sum_in(reg_psum_0_2), .reg_activation(reg_activation_1_2), .reg_weight(reg_weight_1_2), .reg_partial_sum(reg_psum_1_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_3( .activation_in(reg_activation_1_2), .weight_in(reg_weight_0_3), .partial_sum_in(reg_psum_0_3), .reg_activation(reg_activation_1_3), .reg_weight(reg_weight_1_3), .reg_partial_sum(reg_psum_1_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_4( .activation_in(reg_activation_1_3), .weight_in(reg_weight_0_4), .partial_sum_in(reg_psum_0_4), .reg_activation(reg_activation_1_4), .reg_weight(reg_weight_1_4), .reg_partial_sum(reg_psum_1_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_5( .activation_in(reg_activation_1_4), .weight_in(reg_weight_0_5), .partial_sum_in(reg_psum_0_5), .reg_activation(reg_activation_1_5), .reg_weight(reg_weight_1_5), .reg_partial_sum(reg_psum_1_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_6( .activation_in(reg_activation_1_5), .weight_in(reg_weight_0_6), .partial_sum_in(reg_psum_0_6), .reg_activation(reg_activation_1_6), .reg_weight(reg_weight_1_6), .reg_partial_sum(reg_psum_1_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_7( .activation_in(reg_activation_1_6), .weight_in(reg_weight_0_7), .partial_sum_in(reg_psum_0_7), .reg_activation(reg_activation_1_7), .reg_weight(reg_weight_1_7), .reg_partial_sum(reg_psum_1_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_8( .activation_in(reg_activation_1_7), .weight_in(reg_weight_0_8), .partial_sum_in(reg_psum_0_8), .reg_activation(reg_activation_1_8), .reg_weight(reg_weight_1_8), .reg_partial_sum(reg_psum_1_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_9( .activation_in(reg_activation_1_8), .weight_in(reg_weight_0_9), .partial_sum_in(reg_psum_0_9), .reg_activation(reg_activation_1_9), .reg_weight(reg_weight_1_9), .reg_partial_sum(reg_psum_1_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_10( .activation_in(reg_activation_1_9), .weight_in(reg_weight_0_10), .partial_sum_in(reg_psum_0_10), .reg_activation(reg_activation_1_10), .reg_weight(reg_weight_1_10), .reg_partial_sum(reg_psum_1_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_11( .activation_in(reg_activation_1_10), .weight_in(reg_weight_0_11), .partial_sum_in(reg_psum_0_11), .reg_activation(reg_activation_1_11), .reg_weight(reg_weight_1_11), .reg_partial_sum(reg_psum_1_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_12( .activation_in(reg_activation_1_11), .weight_in(reg_weight_0_12), .partial_sum_in(reg_psum_0_12), .reg_activation(reg_activation_1_12), .reg_weight(reg_weight_1_12), .reg_partial_sum(reg_psum_1_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_13( .activation_in(reg_activation_1_12), .weight_in(reg_weight_0_13), .partial_sum_in(reg_psum_0_13), .reg_activation(reg_activation_1_13), .reg_weight(reg_weight_1_13), .reg_partial_sum(reg_psum_1_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_14( .activation_in(reg_activation_1_13), .weight_in(reg_weight_0_14), .partial_sum_in(reg_psum_0_14), .reg_activation(reg_activation_1_14), .reg_weight(reg_weight_1_14), .reg_partial_sum(reg_psum_1_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_15( .activation_in(reg_activation_1_14), .weight_in(reg_weight_0_15), .partial_sum_in(reg_psum_0_15), .reg_activation(reg_activation_1_15), .reg_weight(reg_weight_1_15), .reg_partial_sum(reg_psum_1_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_16( .activation_in(reg_activation_1_15), .weight_in(reg_weight_0_16), .partial_sum_in(reg_psum_0_16), .reg_activation(reg_activation_1_16), .reg_weight(reg_weight_1_16), .reg_partial_sum(reg_psum_1_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_17( .activation_in(reg_activation_1_16), .weight_in(reg_weight_0_17), .partial_sum_in(reg_psum_0_17), .reg_activation(reg_activation_1_17), .reg_weight(reg_weight_1_17), .reg_partial_sum(reg_psum_1_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_18( .activation_in(reg_activation_1_17), .weight_in(reg_weight_0_18), .partial_sum_in(reg_psum_0_18), .reg_activation(reg_activation_1_18), .reg_weight(reg_weight_1_18), .reg_partial_sum(reg_psum_1_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_19( .activation_in(reg_activation_1_18), .weight_in(reg_weight_0_19), .partial_sum_in(reg_psum_0_19), .reg_activation(reg_activation_1_19), .reg_weight(reg_weight_1_19), .reg_partial_sum(reg_psum_1_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_20( .activation_in(reg_activation_1_19), .weight_in(reg_weight_0_20), .partial_sum_in(reg_psum_0_20), .reg_activation(reg_activation_1_20), .reg_weight(reg_weight_1_20), .reg_partial_sum(reg_psum_1_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_21( .activation_in(reg_activation_1_20), .weight_in(reg_weight_0_21), .partial_sum_in(reg_psum_0_21), .reg_activation(reg_activation_1_21), .reg_weight(reg_weight_1_21), .reg_partial_sum(reg_psum_1_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_22( .activation_in(reg_activation_1_21), .weight_in(reg_weight_0_22), .partial_sum_in(reg_psum_0_22), .reg_activation(reg_activation_1_22), .reg_weight(reg_weight_1_22), .reg_partial_sum(reg_psum_1_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_23( .activation_in(reg_activation_1_22), .weight_in(reg_weight_0_23), .partial_sum_in(reg_psum_0_23), .reg_activation(reg_activation_1_23), .reg_weight(reg_weight_1_23), .reg_partial_sum(reg_psum_1_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_24( .activation_in(reg_activation_1_23), .weight_in(reg_weight_0_24), .partial_sum_in(reg_psum_0_24), .reg_activation(reg_activation_1_24), .reg_weight(reg_weight_1_24), .reg_partial_sum(reg_psum_1_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_25( .activation_in(reg_activation_1_24), .weight_in(reg_weight_0_25), .partial_sum_in(reg_psum_0_25), .reg_activation(reg_activation_1_25), .reg_weight(reg_weight_1_25), .reg_partial_sum(reg_psum_1_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_26( .activation_in(reg_activation_1_25), .weight_in(reg_weight_0_26), .partial_sum_in(reg_psum_0_26), .reg_activation(reg_activation_1_26), .reg_weight(reg_weight_1_26), .reg_partial_sum(reg_psum_1_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_27( .activation_in(reg_activation_1_26), .weight_in(reg_weight_0_27), .partial_sum_in(reg_psum_0_27), .reg_activation(reg_activation_1_27), .reg_weight(reg_weight_1_27), .reg_partial_sum(reg_psum_1_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_28( .activation_in(reg_activation_1_27), .weight_in(reg_weight_0_28), .partial_sum_in(reg_psum_0_28), .reg_activation(reg_activation_1_28), .reg_weight(reg_weight_1_28), .reg_partial_sum(reg_psum_1_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_29( .activation_in(reg_activation_1_28), .weight_in(reg_weight_0_29), .partial_sum_in(reg_psum_0_29), .reg_activation(reg_activation_1_29), .reg_weight(reg_weight_1_29), .reg_partial_sum(reg_psum_1_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_30( .activation_in(reg_activation_1_29), .weight_in(reg_weight_0_30), .partial_sum_in(reg_psum_0_30), .reg_activation(reg_activation_1_30), .reg_weight(reg_weight_1_30), .reg_partial_sum(reg_psum_1_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_31( .activation_in(reg_activation_1_30), .weight_in(reg_weight_0_31), .partial_sum_in(reg_psum_0_31), .reg_activation(reg_activation_1_31), .reg_weight(reg_weight_1_31), .reg_partial_sum(reg_psum_1_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_32( .activation_in(reg_activation_1_31), .weight_in(reg_weight_0_32), .partial_sum_in(reg_psum_0_32), .reg_activation(reg_activation_1_32), .reg_weight(reg_weight_1_32), .reg_partial_sum(reg_psum_1_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_33( .activation_in(reg_activation_1_32), .weight_in(reg_weight_0_33), .partial_sum_in(reg_psum_0_33), .reg_activation(reg_activation_1_33), .reg_weight(reg_weight_1_33), .reg_partial_sum(reg_psum_1_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_34( .activation_in(reg_activation_1_33), .weight_in(reg_weight_0_34), .partial_sum_in(reg_psum_0_34), .reg_activation(reg_activation_1_34), .reg_weight(reg_weight_1_34), .reg_partial_sum(reg_psum_1_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_35( .activation_in(reg_activation_1_34), .weight_in(reg_weight_0_35), .partial_sum_in(reg_psum_0_35), .reg_activation(reg_activation_1_35), .reg_weight(reg_weight_1_35), .reg_partial_sum(reg_psum_1_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_36( .activation_in(reg_activation_1_35), .weight_in(reg_weight_0_36), .partial_sum_in(reg_psum_0_36), .reg_activation(reg_activation_1_36), .reg_weight(reg_weight_1_36), .reg_partial_sum(reg_psum_1_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_37( .activation_in(reg_activation_1_36), .weight_in(reg_weight_0_37), .partial_sum_in(reg_psum_0_37), .reg_activation(reg_activation_1_37), .reg_weight(reg_weight_1_37), .reg_partial_sum(reg_psum_1_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_38( .activation_in(reg_activation_1_37), .weight_in(reg_weight_0_38), .partial_sum_in(reg_psum_0_38), .reg_activation(reg_activation_1_38), .reg_weight(reg_weight_1_38), .reg_partial_sum(reg_psum_1_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_39( .activation_in(reg_activation_1_38), .weight_in(reg_weight_0_39), .partial_sum_in(reg_psum_0_39), .reg_activation(reg_activation_1_39), .reg_weight(reg_weight_1_39), .reg_partial_sum(reg_psum_1_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_40( .activation_in(reg_activation_1_39), .weight_in(reg_weight_0_40), .partial_sum_in(reg_psum_0_40), .reg_activation(reg_activation_1_40), .reg_weight(reg_weight_1_40), .reg_partial_sum(reg_psum_1_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_41( .activation_in(reg_activation_1_40), .weight_in(reg_weight_0_41), .partial_sum_in(reg_psum_0_41), .reg_activation(reg_activation_1_41), .reg_weight(reg_weight_1_41), .reg_partial_sum(reg_psum_1_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_42( .activation_in(reg_activation_1_41), .weight_in(reg_weight_0_42), .partial_sum_in(reg_psum_0_42), .reg_activation(reg_activation_1_42), .reg_weight(reg_weight_1_42), .reg_partial_sum(reg_psum_1_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_43( .activation_in(reg_activation_1_42), .weight_in(reg_weight_0_43), .partial_sum_in(reg_psum_0_43), .reg_activation(reg_activation_1_43), .reg_weight(reg_weight_1_43), .reg_partial_sum(reg_psum_1_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_44( .activation_in(reg_activation_1_43), .weight_in(reg_weight_0_44), .partial_sum_in(reg_psum_0_44), .reg_activation(reg_activation_1_44), .reg_weight(reg_weight_1_44), .reg_partial_sum(reg_psum_1_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_45( .activation_in(reg_activation_1_44), .weight_in(reg_weight_0_45), .partial_sum_in(reg_psum_0_45), .reg_activation(reg_activation_1_45), .reg_weight(reg_weight_1_45), .reg_partial_sum(reg_psum_1_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_46( .activation_in(reg_activation_1_45), .weight_in(reg_weight_0_46), .partial_sum_in(reg_psum_0_46), .reg_activation(reg_activation_1_46), .reg_weight(reg_weight_1_46), .reg_partial_sum(reg_psum_1_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_47( .activation_in(reg_activation_1_46), .weight_in(reg_weight_0_47), .partial_sum_in(reg_psum_0_47), .reg_activation(reg_activation_1_47), .reg_weight(reg_weight_1_47), .reg_partial_sum(reg_psum_1_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_48( .activation_in(reg_activation_1_47), .weight_in(reg_weight_0_48), .partial_sum_in(reg_psum_0_48), .reg_activation(reg_activation_1_48), .reg_weight(reg_weight_1_48), .reg_partial_sum(reg_psum_1_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_49( .activation_in(reg_activation_1_48), .weight_in(reg_weight_0_49), .partial_sum_in(reg_psum_0_49), .reg_activation(reg_activation_1_49), .reg_weight(reg_weight_1_49), .reg_partial_sum(reg_psum_1_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_50( .activation_in(reg_activation_1_49), .weight_in(reg_weight_0_50), .partial_sum_in(reg_psum_0_50), .reg_activation(reg_activation_1_50), .reg_weight(reg_weight_1_50), .reg_partial_sum(reg_psum_1_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_51( .activation_in(reg_activation_1_50), .weight_in(reg_weight_0_51), .partial_sum_in(reg_psum_0_51), .reg_activation(reg_activation_1_51), .reg_weight(reg_weight_1_51), .reg_partial_sum(reg_psum_1_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_52( .activation_in(reg_activation_1_51), .weight_in(reg_weight_0_52), .partial_sum_in(reg_psum_0_52), .reg_activation(reg_activation_1_52), .reg_weight(reg_weight_1_52), .reg_partial_sum(reg_psum_1_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_53( .activation_in(reg_activation_1_52), .weight_in(reg_weight_0_53), .partial_sum_in(reg_psum_0_53), .reg_activation(reg_activation_1_53), .reg_weight(reg_weight_1_53), .reg_partial_sum(reg_psum_1_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_54( .activation_in(reg_activation_1_53), .weight_in(reg_weight_0_54), .partial_sum_in(reg_psum_0_54), .reg_activation(reg_activation_1_54), .reg_weight(reg_weight_1_54), .reg_partial_sum(reg_psum_1_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_55( .activation_in(reg_activation_1_54), .weight_in(reg_weight_0_55), .partial_sum_in(reg_psum_0_55), .reg_activation(reg_activation_1_55), .reg_weight(reg_weight_1_55), .reg_partial_sum(reg_psum_1_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_56( .activation_in(reg_activation_1_55), .weight_in(reg_weight_0_56), .partial_sum_in(reg_psum_0_56), .reg_activation(reg_activation_1_56), .reg_weight(reg_weight_1_56), .reg_partial_sum(reg_psum_1_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_57( .activation_in(reg_activation_1_56), .weight_in(reg_weight_0_57), .partial_sum_in(reg_psum_0_57), .reg_activation(reg_activation_1_57), .reg_weight(reg_weight_1_57), .reg_partial_sum(reg_psum_1_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_58( .activation_in(reg_activation_1_57), .weight_in(reg_weight_0_58), .partial_sum_in(reg_psum_0_58), .reg_activation(reg_activation_1_58), .reg_weight(reg_weight_1_58), .reg_partial_sum(reg_psum_1_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_59( .activation_in(reg_activation_1_58), .weight_in(reg_weight_0_59), .partial_sum_in(reg_psum_0_59), .reg_activation(reg_activation_1_59), .reg_weight(reg_weight_1_59), .reg_partial_sum(reg_psum_1_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_60( .activation_in(reg_activation_1_59), .weight_in(reg_weight_0_60), .partial_sum_in(reg_psum_0_60), .reg_activation(reg_activation_1_60), .reg_weight(reg_weight_1_60), .reg_partial_sum(reg_psum_1_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_61( .activation_in(reg_activation_1_60), .weight_in(reg_weight_0_61), .partial_sum_in(reg_psum_0_61), .reg_activation(reg_activation_1_61), .reg_weight(reg_weight_1_61), .reg_partial_sum(reg_psum_1_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_62( .activation_in(reg_activation_1_61), .weight_in(reg_weight_0_62), .partial_sum_in(reg_psum_0_62), .reg_activation(reg_activation_1_62), .reg_weight(reg_weight_1_62), .reg_partial_sum(reg_psum_1_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_63( .activation_in(reg_activation_1_62), .weight_in(reg_weight_0_63), .partial_sum_in(reg_psum_0_63), .reg_weight(reg_weight_1_63), .reg_partial_sum(reg_psum_1_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_0( .activation_in(in_activation_2), .weight_in(reg_weight_1_0), .partial_sum_in(reg_psum_1_0), .reg_activation(reg_activation_2_0), .reg_weight(reg_weight_2_0), .reg_partial_sum(reg_psum_2_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_1( .activation_in(reg_activation_2_0), .weight_in(reg_weight_1_1), .partial_sum_in(reg_psum_1_1), .reg_activation(reg_activation_2_1), .reg_weight(reg_weight_2_1), .reg_partial_sum(reg_psum_2_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_2( .activation_in(reg_activation_2_1), .weight_in(reg_weight_1_2), .partial_sum_in(reg_psum_1_2), .reg_activation(reg_activation_2_2), .reg_weight(reg_weight_2_2), .reg_partial_sum(reg_psum_2_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_3( .activation_in(reg_activation_2_2), .weight_in(reg_weight_1_3), .partial_sum_in(reg_psum_1_3), .reg_activation(reg_activation_2_3), .reg_weight(reg_weight_2_3), .reg_partial_sum(reg_psum_2_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_4( .activation_in(reg_activation_2_3), .weight_in(reg_weight_1_4), .partial_sum_in(reg_psum_1_4), .reg_activation(reg_activation_2_4), .reg_weight(reg_weight_2_4), .reg_partial_sum(reg_psum_2_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_5( .activation_in(reg_activation_2_4), .weight_in(reg_weight_1_5), .partial_sum_in(reg_psum_1_5), .reg_activation(reg_activation_2_5), .reg_weight(reg_weight_2_5), .reg_partial_sum(reg_psum_2_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_6( .activation_in(reg_activation_2_5), .weight_in(reg_weight_1_6), .partial_sum_in(reg_psum_1_6), .reg_activation(reg_activation_2_6), .reg_weight(reg_weight_2_6), .reg_partial_sum(reg_psum_2_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_7( .activation_in(reg_activation_2_6), .weight_in(reg_weight_1_7), .partial_sum_in(reg_psum_1_7), .reg_activation(reg_activation_2_7), .reg_weight(reg_weight_2_7), .reg_partial_sum(reg_psum_2_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_8( .activation_in(reg_activation_2_7), .weight_in(reg_weight_1_8), .partial_sum_in(reg_psum_1_8), .reg_activation(reg_activation_2_8), .reg_weight(reg_weight_2_8), .reg_partial_sum(reg_psum_2_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_9( .activation_in(reg_activation_2_8), .weight_in(reg_weight_1_9), .partial_sum_in(reg_psum_1_9), .reg_activation(reg_activation_2_9), .reg_weight(reg_weight_2_9), .reg_partial_sum(reg_psum_2_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_10( .activation_in(reg_activation_2_9), .weight_in(reg_weight_1_10), .partial_sum_in(reg_psum_1_10), .reg_activation(reg_activation_2_10), .reg_weight(reg_weight_2_10), .reg_partial_sum(reg_psum_2_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_11( .activation_in(reg_activation_2_10), .weight_in(reg_weight_1_11), .partial_sum_in(reg_psum_1_11), .reg_activation(reg_activation_2_11), .reg_weight(reg_weight_2_11), .reg_partial_sum(reg_psum_2_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_12( .activation_in(reg_activation_2_11), .weight_in(reg_weight_1_12), .partial_sum_in(reg_psum_1_12), .reg_activation(reg_activation_2_12), .reg_weight(reg_weight_2_12), .reg_partial_sum(reg_psum_2_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_13( .activation_in(reg_activation_2_12), .weight_in(reg_weight_1_13), .partial_sum_in(reg_psum_1_13), .reg_activation(reg_activation_2_13), .reg_weight(reg_weight_2_13), .reg_partial_sum(reg_psum_2_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_14( .activation_in(reg_activation_2_13), .weight_in(reg_weight_1_14), .partial_sum_in(reg_psum_1_14), .reg_activation(reg_activation_2_14), .reg_weight(reg_weight_2_14), .reg_partial_sum(reg_psum_2_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_15( .activation_in(reg_activation_2_14), .weight_in(reg_weight_1_15), .partial_sum_in(reg_psum_1_15), .reg_activation(reg_activation_2_15), .reg_weight(reg_weight_2_15), .reg_partial_sum(reg_psum_2_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_16( .activation_in(reg_activation_2_15), .weight_in(reg_weight_1_16), .partial_sum_in(reg_psum_1_16), .reg_activation(reg_activation_2_16), .reg_weight(reg_weight_2_16), .reg_partial_sum(reg_psum_2_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_17( .activation_in(reg_activation_2_16), .weight_in(reg_weight_1_17), .partial_sum_in(reg_psum_1_17), .reg_activation(reg_activation_2_17), .reg_weight(reg_weight_2_17), .reg_partial_sum(reg_psum_2_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_18( .activation_in(reg_activation_2_17), .weight_in(reg_weight_1_18), .partial_sum_in(reg_psum_1_18), .reg_activation(reg_activation_2_18), .reg_weight(reg_weight_2_18), .reg_partial_sum(reg_psum_2_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_19( .activation_in(reg_activation_2_18), .weight_in(reg_weight_1_19), .partial_sum_in(reg_psum_1_19), .reg_activation(reg_activation_2_19), .reg_weight(reg_weight_2_19), .reg_partial_sum(reg_psum_2_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_20( .activation_in(reg_activation_2_19), .weight_in(reg_weight_1_20), .partial_sum_in(reg_psum_1_20), .reg_activation(reg_activation_2_20), .reg_weight(reg_weight_2_20), .reg_partial_sum(reg_psum_2_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_21( .activation_in(reg_activation_2_20), .weight_in(reg_weight_1_21), .partial_sum_in(reg_psum_1_21), .reg_activation(reg_activation_2_21), .reg_weight(reg_weight_2_21), .reg_partial_sum(reg_psum_2_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_22( .activation_in(reg_activation_2_21), .weight_in(reg_weight_1_22), .partial_sum_in(reg_psum_1_22), .reg_activation(reg_activation_2_22), .reg_weight(reg_weight_2_22), .reg_partial_sum(reg_psum_2_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_23( .activation_in(reg_activation_2_22), .weight_in(reg_weight_1_23), .partial_sum_in(reg_psum_1_23), .reg_activation(reg_activation_2_23), .reg_weight(reg_weight_2_23), .reg_partial_sum(reg_psum_2_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_24( .activation_in(reg_activation_2_23), .weight_in(reg_weight_1_24), .partial_sum_in(reg_psum_1_24), .reg_activation(reg_activation_2_24), .reg_weight(reg_weight_2_24), .reg_partial_sum(reg_psum_2_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_25( .activation_in(reg_activation_2_24), .weight_in(reg_weight_1_25), .partial_sum_in(reg_psum_1_25), .reg_activation(reg_activation_2_25), .reg_weight(reg_weight_2_25), .reg_partial_sum(reg_psum_2_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_26( .activation_in(reg_activation_2_25), .weight_in(reg_weight_1_26), .partial_sum_in(reg_psum_1_26), .reg_activation(reg_activation_2_26), .reg_weight(reg_weight_2_26), .reg_partial_sum(reg_psum_2_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_27( .activation_in(reg_activation_2_26), .weight_in(reg_weight_1_27), .partial_sum_in(reg_psum_1_27), .reg_activation(reg_activation_2_27), .reg_weight(reg_weight_2_27), .reg_partial_sum(reg_psum_2_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_28( .activation_in(reg_activation_2_27), .weight_in(reg_weight_1_28), .partial_sum_in(reg_psum_1_28), .reg_activation(reg_activation_2_28), .reg_weight(reg_weight_2_28), .reg_partial_sum(reg_psum_2_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_29( .activation_in(reg_activation_2_28), .weight_in(reg_weight_1_29), .partial_sum_in(reg_psum_1_29), .reg_activation(reg_activation_2_29), .reg_weight(reg_weight_2_29), .reg_partial_sum(reg_psum_2_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_30( .activation_in(reg_activation_2_29), .weight_in(reg_weight_1_30), .partial_sum_in(reg_psum_1_30), .reg_activation(reg_activation_2_30), .reg_weight(reg_weight_2_30), .reg_partial_sum(reg_psum_2_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_31( .activation_in(reg_activation_2_30), .weight_in(reg_weight_1_31), .partial_sum_in(reg_psum_1_31), .reg_activation(reg_activation_2_31), .reg_weight(reg_weight_2_31), .reg_partial_sum(reg_psum_2_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_32( .activation_in(reg_activation_2_31), .weight_in(reg_weight_1_32), .partial_sum_in(reg_psum_1_32), .reg_activation(reg_activation_2_32), .reg_weight(reg_weight_2_32), .reg_partial_sum(reg_psum_2_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_33( .activation_in(reg_activation_2_32), .weight_in(reg_weight_1_33), .partial_sum_in(reg_psum_1_33), .reg_activation(reg_activation_2_33), .reg_weight(reg_weight_2_33), .reg_partial_sum(reg_psum_2_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_34( .activation_in(reg_activation_2_33), .weight_in(reg_weight_1_34), .partial_sum_in(reg_psum_1_34), .reg_activation(reg_activation_2_34), .reg_weight(reg_weight_2_34), .reg_partial_sum(reg_psum_2_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_35( .activation_in(reg_activation_2_34), .weight_in(reg_weight_1_35), .partial_sum_in(reg_psum_1_35), .reg_activation(reg_activation_2_35), .reg_weight(reg_weight_2_35), .reg_partial_sum(reg_psum_2_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_36( .activation_in(reg_activation_2_35), .weight_in(reg_weight_1_36), .partial_sum_in(reg_psum_1_36), .reg_activation(reg_activation_2_36), .reg_weight(reg_weight_2_36), .reg_partial_sum(reg_psum_2_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_37( .activation_in(reg_activation_2_36), .weight_in(reg_weight_1_37), .partial_sum_in(reg_psum_1_37), .reg_activation(reg_activation_2_37), .reg_weight(reg_weight_2_37), .reg_partial_sum(reg_psum_2_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_38( .activation_in(reg_activation_2_37), .weight_in(reg_weight_1_38), .partial_sum_in(reg_psum_1_38), .reg_activation(reg_activation_2_38), .reg_weight(reg_weight_2_38), .reg_partial_sum(reg_psum_2_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_39( .activation_in(reg_activation_2_38), .weight_in(reg_weight_1_39), .partial_sum_in(reg_psum_1_39), .reg_activation(reg_activation_2_39), .reg_weight(reg_weight_2_39), .reg_partial_sum(reg_psum_2_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_40( .activation_in(reg_activation_2_39), .weight_in(reg_weight_1_40), .partial_sum_in(reg_psum_1_40), .reg_activation(reg_activation_2_40), .reg_weight(reg_weight_2_40), .reg_partial_sum(reg_psum_2_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_41( .activation_in(reg_activation_2_40), .weight_in(reg_weight_1_41), .partial_sum_in(reg_psum_1_41), .reg_activation(reg_activation_2_41), .reg_weight(reg_weight_2_41), .reg_partial_sum(reg_psum_2_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_42( .activation_in(reg_activation_2_41), .weight_in(reg_weight_1_42), .partial_sum_in(reg_psum_1_42), .reg_activation(reg_activation_2_42), .reg_weight(reg_weight_2_42), .reg_partial_sum(reg_psum_2_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_43( .activation_in(reg_activation_2_42), .weight_in(reg_weight_1_43), .partial_sum_in(reg_psum_1_43), .reg_activation(reg_activation_2_43), .reg_weight(reg_weight_2_43), .reg_partial_sum(reg_psum_2_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_44( .activation_in(reg_activation_2_43), .weight_in(reg_weight_1_44), .partial_sum_in(reg_psum_1_44), .reg_activation(reg_activation_2_44), .reg_weight(reg_weight_2_44), .reg_partial_sum(reg_psum_2_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_45( .activation_in(reg_activation_2_44), .weight_in(reg_weight_1_45), .partial_sum_in(reg_psum_1_45), .reg_activation(reg_activation_2_45), .reg_weight(reg_weight_2_45), .reg_partial_sum(reg_psum_2_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_46( .activation_in(reg_activation_2_45), .weight_in(reg_weight_1_46), .partial_sum_in(reg_psum_1_46), .reg_activation(reg_activation_2_46), .reg_weight(reg_weight_2_46), .reg_partial_sum(reg_psum_2_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_47( .activation_in(reg_activation_2_46), .weight_in(reg_weight_1_47), .partial_sum_in(reg_psum_1_47), .reg_activation(reg_activation_2_47), .reg_weight(reg_weight_2_47), .reg_partial_sum(reg_psum_2_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_48( .activation_in(reg_activation_2_47), .weight_in(reg_weight_1_48), .partial_sum_in(reg_psum_1_48), .reg_activation(reg_activation_2_48), .reg_weight(reg_weight_2_48), .reg_partial_sum(reg_psum_2_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_49( .activation_in(reg_activation_2_48), .weight_in(reg_weight_1_49), .partial_sum_in(reg_psum_1_49), .reg_activation(reg_activation_2_49), .reg_weight(reg_weight_2_49), .reg_partial_sum(reg_psum_2_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_50( .activation_in(reg_activation_2_49), .weight_in(reg_weight_1_50), .partial_sum_in(reg_psum_1_50), .reg_activation(reg_activation_2_50), .reg_weight(reg_weight_2_50), .reg_partial_sum(reg_psum_2_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_51( .activation_in(reg_activation_2_50), .weight_in(reg_weight_1_51), .partial_sum_in(reg_psum_1_51), .reg_activation(reg_activation_2_51), .reg_weight(reg_weight_2_51), .reg_partial_sum(reg_psum_2_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_52( .activation_in(reg_activation_2_51), .weight_in(reg_weight_1_52), .partial_sum_in(reg_psum_1_52), .reg_activation(reg_activation_2_52), .reg_weight(reg_weight_2_52), .reg_partial_sum(reg_psum_2_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_53( .activation_in(reg_activation_2_52), .weight_in(reg_weight_1_53), .partial_sum_in(reg_psum_1_53), .reg_activation(reg_activation_2_53), .reg_weight(reg_weight_2_53), .reg_partial_sum(reg_psum_2_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_54( .activation_in(reg_activation_2_53), .weight_in(reg_weight_1_54), .partial_sum_in(reg_psum_1_54), .reg_activation(reg_activation_2_54), .reg_weight(reg_weight_2_54), .reg_partial_sum(reg_psum_2_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_55( .activation_in(reg_activation_2_54), .weight_in(reg_weight_1_55), .partial_sum_in(reg_psum_1_55), .reg_activation(reg_activation_2_55), .reg_weight(reg_weight_2_55), .reg_partial_sum(reg_psum_2_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_56( .activation_in(reg_activation_2_55), .weight_in(reg_weight_1_56), .partial_sum_in(reg_psum_1_56), .reg_activation(reg_activation_2_56), .reg_weight(reg_weight_2_56), .reg_partial_sum(reg_psum_2_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_57( .activation_in(reg_activation_2_56), .weight_in(reg_weight_1_57), .partial_sum_in(reg_psum_1_57), .reg_activation(reg_activation_2_57), .reg_weight(reg_weight_2_57), .reg_partial_sum(reg_psum_2_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_58( .activation_in(reg_activation_2_57), .weight_in(reg_weight_1_58), .partial_sum_in(reg_psum_1_58), .reg_activation(reg_activation_2_58), .reg_weight(reg_weight_2_58), .reg_partial_sum(reg_psum_2_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_59( .activation_in(reg_activation_2_58), .weight_in(reg_weight_1_59), .partial_sum_in(reg_psum_1_59), .reg_activation(reg_activation_2_59), .reg_weight(reg_weight_2_59), .reg_partial_sum(reg_psum_2_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_60( .activation_in(reg_activation_2_59), .weight_in(reg_weight_1_60), .partial_sum_in(reg_psum_1_60), .reg_activation(reg_activation_2_60), .reg_weight(reg_weight_2_60), .reg_partial_sum(reg_psum_2_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_61( .activation_in(reg_activation_2_60), .weight_in(reg_weight_1_61), .partial_sum_in(reg_psum_1_61), .reg_activation(reg_activation_2_61), .reg_weight(reg_weight_2_61), .reg_partial_sum(reg_psum_2_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_62( .activation_in(reg_activation_2_61), .weight_in(reg_weight_1_62), .partial_sum_in(reg_psum_1_62), .reg_activation(reg_activation_2_62), .reg_weight(reg_weight_2_62), .reg_partial_sum(reg_psum_2_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_63( .activation_in(reg_activation_2_62), .weight_in(reg_weight_1_63), .partial_sum_in(reg_psum_1_63), .reg_weight(reg_weight_2_63), .reg_partial_sum(reg_psum_2_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_0( .activation_in(in_activation_3), .weight_in(reg_weight_2_0), .partial_sum_in(reg_psum_2_0), .reg_activation(reg_activation_3_0), .reg_weight(reg_weight_3_0), .reg_partial_sum(reg_psum_3_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_1( .activation_in(reg_activation_3_0), .weight_in(reg_weight_2_1), .partial_sum_in(reg_psum_2_1), .reg_activation(reg_activation_3_1), .reg_weight(reg_weight_3_1), .reg_partial_sum(reg_psum_3_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_2( .activation_in(reg_activation_3_1), .weight_in(reg_weight_2_2), .partial_sum_in(reg_psum_2_2), .reg_activation(reg_activation_3_2), .reg_weight(reg_weight_3_2), .reg_partial_sum(reg_psum_3_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_3( .activation_in(reg_activation_3_2), .weight_in(reg_weight_2_3), .partial_sum_in(reg_psum_2_3), .reg_activation(reg_activation_3_3), .reg_weight(reg_weight_3_3), .reg_partial_sum(reg_psum_3_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_4( .activation_in(reg_activation_3_3), .weight_in(reg_weight_2_4), .partial_sum_in(reg_psum_2_4), .reg_activation(reg_activation_3_4), .reg_weight(reg_weight_3_4), .reg_partial_sum(reg_psum_3_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_5( .activation_in(reg_activation_3_4), .weight_in(reg_weight_2_5), .partial_sum_in(reg_psum_2_5), .reg_activation(reg_activation_3_5), .reg_weight(reg_weight_3_5), .reg_partial_sum(reg_psum_3_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_6( .activation_in(reg_activation_3_5), .weight_in(reg_weight_2_6), .partial_sum_in(reg_psum_2_6), .reg_activation(reg_activation_3_6), .reg_weight(reg_weight_3_6), .reg_partial_sum(reg_psum_3_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_7( .activation_in(reg_activation_3_6), .weight_in(reg_weight_2_7), .partial_sum_in(reg_psum_2_7), .reg_activation(reg_activation_3_7), .reg_weight(reg_weight_3_7), .reg_partial_sum(reg_psum_3_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_8( .activation_in(reg_activation_3_7), .weight_in(reg_weight_2_8), .partial_sum_in(reg_psum_2_8), .reg_activation(reg_activation_3_8), .reg_weight(reg_weight_3_8), .reg_partial_sum(reg_psum_3_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_9( .activation_in(reg_activation_3_8), .weight_in(reg_weight_2_9), .partial_sum_in(reg_psum_2_9), .reg_activation(reg_activation_3_9), .reg_weight(reg_weight_3_9), .reg_partial_sum(reg_psum_3_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_10( .activation_in(reg_activation_3_9), .weight_in(reg_weight_2_10), .partial_sum_in(reg_psum_2_10), .reg_activation(reg_activation_3_10), .reg_weight(reg_weight_3_10), .reg_partial_sum(reg_psum_3_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_11( .activation_in(reg_activation_3_10), .weight_in(reg_weight_2_11), .partial_sum_in(reg_psum_2_11), .reg_activation(reg_activation_3_11), .reg_weight(reg_weight_3_11), .reg_partial_sum(reg_psum_3_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_12( .activation_in(reg_activation_3_11), .weight_in(reg_weight_2_12), .partial_sum_in(reg_psum_2_12), .reg_activation(reg_activation_3_12), .reg_weight(reg_weight_3_12), .reg_partial_sum(reg_psum_3_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_13( .activation_in(reg_activation_3_12), .weight_in(reg_weight_2_13), .partial_sum_in(reg_psum_2_13), .reg_activation(reg_activation_3_13), .reg_weight(reg_weight_3_13), .reg_partial_sum(reg_psum_3_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_14( .activation_in(reg_activation_3_13), .weight_in(reg_weight_2_14), .partial_sum_in(reg_psum_2_14), .reg_activation(reg_activation_3_14), .reg_weight(reg_weight_3_14), .reg_partial_sum(reg_psum_3_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_15( .activation_in(reg_activation_3_14), .weight_in(reg_weight_2_15), .partial_sum_in(reg_psum_2_15), .reg_activation(reg_activation_3_15), .reg_weight(reg_weight_3_15), .reg_partial_sum(reg_psum_3_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_16( .activation_in(reg_activation_3_15), .weight_in(reg_weight_2_16), .partial_sum_in(reg_psum_2_16), .reg_activation(reg_activation_3_16), .reg_weight(reg_weight_3_16), .reg_partial_sum(reg_psum_3_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_17( .activation_in(reg_activation_3_16), .weight_in(reg_weight_2_17), .partial_sum_in(reg_psum_2_17), .reg_activation(reg_activation_3_17), .reg_weight(reg_weight_3_17), .reg_partial_sum(reg_psum_3_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_18( .activation_in(reg_activation_3_17), .weight_in(reg_weight_2_18), .partial_sum_in(reg_psum_2_18), .reg_activation(reg_activation_3_18), .reg_weight(reg_weight_3_18), .reg_partial_sum(reg_psum_3_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_19( .activation_in(reg_activation_3_18), .weight_in(reg_weight_2_19), .partial_sum_in(reg_psum_2_19), .reg_activation(reg_activation_3_19), .reg_weight(reg_weight_3_19), .reg_partial_sum(reg_psum_3_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_20( .activation_in(reg_activation_3_19), .weight_in(reg_weight_2_20), .partial_sum_in(reg_psum_2_20), .reg_activation(reg_activation_3_20), .reg_weight(reg_weight_3_20), .reg_partial_sum(reg_psum_3_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_21( .activation_in(reg_activation_3_20), .weight_in(reg_weight_2_21), .partial_sum_in(reg_psum_2_21), .reg_activation(reg_activation_3_21), .reg_weight(reg_weight_3_21), .reg_partial_sum(reg_psum_3_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_22( .activation_in(reg_activation_3_21), .weight_in(reg_weight_2_22), .partial_sum_in(reg_psum_2_22), .reg_activation(reg_activation_3_22), .reg_weight(reg_weight_3_22), .reg_partial_sum(reg_psum_3_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_23( .activation_in(reg_activation_3_22), .weight_in(reg_weight_2_23), .partial_sum_in(reg_psum_2_23), .reg_activation(reg_activation_3_23), .reg_weight(reg_weight_3_23), .reg_partial_sum(reg_psum_3_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_24( .activation_in(reg_activation_3_23), .weight_in(reg_weight_2_24), .partial_sum_in(reg_psum_2_24), .reg_activation(reg_activation_3_24), .reg_weight(reg_weight_3_24), .reg_partial_sum(reg_psum_3_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_25( .activation_in(reg_activation_3_24), .weight_in(reg_weight_2_25), .partial_sum_in(reg_psum_2_25), .reg_activation(reg_activation_3_25), .reg_weight(reg_weight_3_25), .reg_partial_sum(reg_psum_3_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_26( .activation_in(reg_activation_3_25), .weight_in(reg_weight_2_26), .partial_sum_in(reg_psum_2_26), .reg_activation(reg_activation_3_26), .reg_weight(reg_weight_3_26), .reg_partial_sum(reg_psum_3_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_27( .activation_in(reg_activation_3_26), .weight_in(reg_weight_2_27), .partial_sum_in(reg_psum_2_27), .reg_activation(reg_activation_3_27), .reg_weight(reg_weight_3_27), .reg_partial_sum(reg_psum_3_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_28( .activation_in(reg_activation_3_27), .weight_in(reg_weight_2_28), .partial_sum_in(reg_psum_2_28), .reg_activation(reg_activation_3_28), .reg_weight(reg_weight_3_28), .reg_partial_sum(reg_psum_3_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_29( .activation_in(reg_activation_3_28), .weight_in(reg_weight_2_29), .partial_sum_in(reg_psum_2_29), .reg_activation(reg_activation_3_29), .reg_weight(reg_weight_3_29), .reg_partial_sum(reg_psum_3_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_30( .activation_in(reg_activation_3_29), .weight_in(reg_weight_2_30), .partial_sum_in(reg_psum_2_30), .reg_activation(reg_activation_3_30), .reg_weight(reg_weight_3_30), .reg_partial_sum(reg_psum_3_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_31( .activation_in(reg_activation_3_30), .weight_in(reg_weight_2_31), .partial_sum_in(reg_psum_2_31), .reg_activation(reg_activation_3_31), .reg_weight(reg_weight_3_31), .reg_partial_sum(reg_psum_3_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_32( .activation_in(reg_activation_3_31), .weight_in(reg_weight_2_32), .partial_sum_in(reg_psum_2_32), .reg_activation(reg_activation_3_32), .reg_weight(reg_weight_3_32), .reg_partial_sum(reg_psum_3_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_33( .activation_in(reg_activation_3_32), .weight_in(reg_weight_2_33), .partial_sum_in(reg_psum_2_33), .reg_activation(reg_activation_3_33), .reg_weight(reg_weight_3_33), .reg_partial_sum(reg_psum_3_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_34( .activation_in(reg_activation_3_33), .weight_in(reg_weight_2_34), .partial_sum_in(reg_psum_2_34), .reg_activation(reg_activation_3_34), .reg_weight(reg_weight_3_34), .reg_partial_sum(reg_psum_3_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_35( .activation_in(reg_activation_3_34), .weight_in(reg_weight_2_35), .partial_sum_in(reg_psum_2_35), .reg_activation(reg_activation_3_35), .reg_weight(reg_weight_3_35), .reg_partial_sum(reg_psum_3_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_36( .activation_in(reg_activation_3_35), .weight_in(reg_weight_2_36), .partial_sum_in(reg_psum_2_36), .reg_activation(reg_activation_3_36), .reg_weight(reg_weight_3_36), .reg_partial_sum(reg_psum_3_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_37( .activation_in(reg_activation_3_36), .weight_in(reg_weight_2_37), .partial_sum_in(reg_psum_2_37), .reg_activation(reg_activation_3_37), .reg_weight(reg_weight_3_37), .reg_partial_sum(reg_psum_3_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_38( .activation_in(reg_activation_3_37), .weight_in(reg_weight_2_38), .partial_sum_in(reg_psum_2_38), .reg_activation(reg_activation_3_38), .reg_weight(reg_weight_3_38), .reg_partial_sum(reg_psum_3_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_39( .activation_in(reg_activation_3_38), .weight_in(reg_weight_2_39), .partial_sum_in(reg_psum_2_39), .reg_activation(reg_activation_3_39), .reg_weight(reg_weight_3_39), .reg_partial_sum(reg_psum_3_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_40( .activation_in(reg_activation_3_39), .weight_in(reg_weight_2_40), .partial_sum_in(reg_psum_2_40), .reg_activation(reg_activation_3_40), .reg_weight(reg_weight_3_40), .reg_partial_sum(reg_psum_3_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_41( .activation_in(reg_activation_3_40), .weight_in(reg_weight_2_41), .partial_sum_in(reg_psum_2_41), .reg_activation(reg_activation_3_41), .reg_weight(reg_weight_3_41), .reg_partial_sum(reg_psum_3_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_42( .activation_in(reg_activation_3_41), .weight_in(reg_weight_2_42), .partial_sum_in(reg_psum_2_42), .reg_activation(reg_activation_3_42), .reg_weight(reg_weight_3_42), .reg_partial_sum(reg_psum_3_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_43( .activation_in(reg_activation_3_42), .weight_in(reg_weight_2_43), .partial_sum_in(reg_psum_2_43), .reg_activation(reg_activation_3_43), .reg_weight(reg_weight_3_43), .reg_partial_sum(reg_psum_3_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_44( .activation_in(reg_activation_3_43), .weight_in(reg_weight_2_44), .partial_sum_in(reg_psum_2_44), .reg_activation(reg_activation_3_44), .reg_weight(reg_weight_3_44), .reg_partial_sum(reg_psum_3_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_45( .activation_in(reg_activation_3_44), .weight_in(reg_weight_2_45), .partial_sum_in(reg_psum_2_45), .reg_activation(reg_activation_3_45), .reg_weight(reg_weight_3_45), .reg_partial_sum(reg_psum_3_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_46( .activation_in(reg_activation_3_45), .weight_in(reg_weight_2_46), .partial_sum_in(reg_psum_2_46), .reg_activation(reg_activation_3_46), .reg_weight(reg_weight_3_46), .reg_partial_sum(reg_psum_3_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_47( .activation_in(reg_activation_3_46), .weight_in(reg_weight_2_47), .partial_sum_in(reg_psum_2_47), .reg_activation(reg_activation_3_47), .reg_weight(reg_weight_3_47), .reg_partial_sum(reg_psum_3_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_48( .activation_in(reg_activation_3_47), .weight_in(reg_weight_2_48), .partial_sum_in(reg_psum_2_48), .reg_activation(reg_activation_3_48), .reg_weight(reg_weight_3_48), .reg_partial_sum(reg_psum_3_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_49( .activation_in(reg_activation_3_48), .weight_in(reg_weight_2_49), .partial_sum_in(reg_psum_2_49), .reg_activation(reg_activation_3_49), .reg_weight(reg_weight_3_49), .reg_partial_sum(reg_psum_3_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_50( .activation_in(reg_activation_3_49), .weight_in(reg_weight_2_50), .partial_sum_in(reg_psum_2_50), .reg_activation(reg_activation_3_50), .reg_weight(reg_weight_3_50), .reg_partial_sum(reg_psum_3_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_51( .activation_in(reg_activation_3_50), .weight_in(reg_weight_2_51), .partial_sum_in(reg_psum_2_51), .reg_activation(reg_activation_3_51), .reg_weight(reg_weight_3_51), .reg_partial_sum(reg_psum_3_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_52( .activation_in(reg_activation_3_51), .weight_in(reg_weight_2_52), .partial_sum_in(reg_psum_2_52), .reg_activation(reg_activation_3_52), .reg_weight(reg_weight_3_52), .reg_partial_sum(reg_psum_3_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_53( .activation_in(reg_activation_3_52), .weight_in(reg_weight_2_53), .partial_sum_in(reg_psum_2_53), .reg_activation(reg_activation_3_53), .reg_weight(reg_weight_3_53), .reg_partial_sum(reg_psum_3_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_54( .activation_in(reg_activation_3_53), .weight_in(reg_weight_2_54), .partial_sum_in(reg_psum_2_54), .reg_activation(reg_activation_3_54), .reg_weight(reg_weight_3_54), .reg_partial_sum(reg_psum_3_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_55( .activation_in(reg_activation_3_54), .weight_in(reg_weight_2_55), .partial_sum_in(reg_psum_2_55), .reg_activation(reg_activation_3_55), .reg_weight(reg_weight_3_55), .reg_partial_sum(reg_psum_3_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_56( .activation_in(reg_activation_3_55), .weight_in(reg_weight_2_56), .partial_sum_in(reg_psum_2_56), .reg_activation(reg_activation_3_56), .reg_weight(reg_weight_3_56), .reg_partial_sum(reg_psum_3_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_57( .activation_in(reg_activation_3_56), .weight_in(reg_weight_2_57), .partial_sum_in(reg_psum_2_57), .reg_activation(reg_activation_3_57), .reg_weight(reg_weight_3_57), .reg_partial_sum(reg_psum_3_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_58( .activation_in(reg_activation_3_57), .weight_in(reg_weight_2_58), .partial_sum_in(reg_psum_2_58), .reg_activation(reg_activation_3_58), .reg_weight(reg_weight_3_58), .reg_partial_sum(reg_psum_3_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_59( .activation_in(reg_activation_3_58), .weight_in(reg_weight_2_59), .partial_sum_in(reg_psum_2_59), .reg_activation(reg_activation_3_59), .reg_weight(reg_weight_3_59), .reg_partial_sum(reg_psum_3_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_60( .activation_in(reg_activation_3_59), .weight_in(reg_weight_2_60), .partial_sum_in(reg_psum_2_60), .reg_activation(reg_activation_3_60), .reg_weight(reg_weight_3_60), .reg_partial_sum(reg_psum_3_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_61( .activation_in(reg_activation_3_60), .weight_in(reg_weight_2_61), .partial_sum_in(reg_psum_2_61), .reg_activation(reg_activation_3_61), .reg_weight(reg_weight_3_61), .reg_partial_sum(reg_psum_3_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_62( .activation_in(reg_activation_3_61), .weight_in(reg_weight_2_62), .partial_sum_in(reg_psum_2_62), .reg_activation(reg_activation_3_62), .reg_weight(reg_weight_3_62), .reg_partial_sum(reg_psum_3_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_63( .activation_in(reg_activation_3_62), .weight_in(reg_weight_2_63), .partial_sum_in(reg_psum_2_63), .reg_weight(reg_weight_3_63), .reg_partial_sum(reg_psum_3_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_0( .activation_in(in_activation_4), .weight_in(reg_weight_3_0), .partial_sum_in(reg_psum_3_0), .reg_activation(reg_activation_4_0), .reg_weight(reg_weight_4_0), .reg_partial_sum(reg_psum_4_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_1( .activation_in(reg_activation_4_0), .weight_in(reg_weight_3_1), .partial_sum_in(reg_psum_3_1), .reg_activation(reg_activation_4_1), .reg_weight(reg_weight_4_1), .reg_partial_sum(reg_psum_4_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_2( .activation_in(reg_activation_4_1), .weight_in(reg_weight_3_2), .partial_sum_in(reg_psum_3_2), .reg_activation(reg_activation_4_2), .reg_weight(reg_weight_4_2), .reg_partial_sum(reg_psum_4_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_3( .activation_in(reg_activation_4_2), .weight_in(reg_weight_3_3), .partial_sum_in(reg_psum_3_3), .reg_activation(reg_activation_4_3), .reg_weight(reg_weight_4_3), .reg_partial_sum(reg_psum_4_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_4( .activation_in(reg_activation_4_3), .weight_in(reg_weight_3_4), .partial_sum_in(reg_psum_3_4), .reg_activation(reg_activation_4_4), .reg_weight(reg_weight_4_4), .reg_partial_sum(reg_psum_4_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_5( .activation_in(reg_activation_4_4), .weight_in(reg_weight_3_5), .partial_sum_in(reg_psum_3_5), .reg_activation(reg_activation_4_5), .reg_weight(reg_weight_4_5), .reg_partial_sum(reg_psum_4_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_6( .activation_in(reg_activation_4_5), .weight_in(reg_weight_3_6), .partial_sum_in(reg_psum_3_6), .reg_activation(reg_activation_4_6), .reg_weight(reg_weight_4_6), .reg_partial_sum(reg_psum_4_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_7( .activation_in(reg_activation_4_6), .weight_in(reg_weight_3_7), .partial_sum_in(reg_psum_3_7), .reg_activation(reg_activation_4_7), .reg_weight(reg_weight_4_7), .reg_partial_sum(reg_psum_4_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_8( .activation_in(reg_activation_4_7), .weight_in(reg_weight_3_8), .partial_sum_in(reg_psum_3_8), .reg_activation(reg_activation_4_8), .reg_weight(reg_weight_4_8), .reg_partial_sum(reg_psum_4_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_9( .activation_in(reg_activation_4_8), .weight_in(reg_weight_3_9), .partial_sum_in(reg_psum_3_9), .reg_activation(reg_activation_4_9), .reg_weight(reg_weight_4_9), .reg_partial_sum(reg_psum_4_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_10( .activation_in(reg_activation_4_9), .weight_in(reg_weight_3_10), .partial_sum_in(reg_psum_3_10), .reg_activation(reg_activation_4_10), .reg_weight(reg_weight_4_10), .reg_partial_sum(reg_psum_4_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_11( .activation_in(reg_activation_4_10), .weight_in(reg_weight_3_11), .partial_sum_in(reg_psum_3_11), .reg_activation(reg_activation_4_11), .reg_weight(reg_weight_4_11), .reg_partial_sum(reg_psum_4_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_12( .activation_in(reg_activation_4_11), .weight_in(reg_weight_3_12), .partial_sum_in(reg_psum_3_12), .reg_activation(reg_activation_4_12), .reg_weight(reg_weight_4_12), .reg_partial_sum(reg_psum_4_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_13( .activation_in(reg_activation_4_12), .weight_in(reg_weight_3_13), .partial_sum_in(reg_psum_3_13), .reg_activation(reg_activation_4_13), .reg_weight(reg_weight_4_13), .reg_partial_sum(reg_psum_4_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_14( .activation_in(reg_activation_4_13), .weight_in(reg_weight_3_14), .partial_sum_in(reg_psum_3_14), .reg_activation(reg_activation_4_14), .reg_weight(reg_weight_4_14), .reg_partial_sum(reg_psum_4_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_15( .activation_in(reg_activation_4_14), .weight_in(reg_weight_3_15), .partial_sum_in(reg_psum_3_15), .reg_activation(reg_activation_4_15), .reg_weight(reg_weight_4_15), .reg_partial_sum(reg_psum_4_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_16( .activation_in(reg_activation_4_15), .weight_in(reg_weight_3_16), .partial_sum_in(reg_psum_3_16), .reg_activation(reg_activation_4_16), .reg_weight(reg_weight_4_16), .reg_partial_sum(reg_psum_4_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_17( .activation_in(reg_activation_4_16), .weight_in(reg_weight_3_17), .partial_sum_in(reg_psum_3_17), .reg_activation(reg_activation_4_17), .reg_weight(reg_weight_4_17), .reg_partial_sum(reg_psum_4_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_18( .activation_in(reg_activation_4_17), .weight_in(reg_weight_3_18), .partial_sum_in(reg_psum_3_18), .reg_activation(reg_activation_4_18), .reg_weight(reg_weight_4_18), .reg_partial_sum(reg_psum_4_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_19( .activation_in(reg_activation_4_18), .weight_in(reg_weight_3_19), .partial_sum_in(reg_psum_3_19), .reg_activation(reg_activation_4_19), .reg_weight(reg_weight_4_19), .reg_partial_sum(reg_psum_4_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_20( .activation_in(reg_activation_4_19), .weight_in(reg_weight_3_20), .partial_sum_in(reg_psum_3_20), .reg_activation(reg_activation_4_20), .reg_weight(reg_weight_4_20), .reg_partial_sum(reg_psum_4_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_21( .activation_in(reg_activation_4_20), .weight_in(reg_weight_3_21), .partial_sum_in(reg_psum_3_21), .reg_activation(reg_activation_4_21), .reg_weight(reg_weight_4_21), .reg_partial_sum(reg_psum_4_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_22( .activation_in(reg_activation_4_21), .weight_in(reg_weight_3_22), .partial_sum_in(reg_psum_3_22), .reg_activation(reg_activation_4_22), .reg_weight(reg_weight_4_22), .reg_partial_sum(reg_psum_4_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_23( .activation_in(reg_activation_4_22), .weight_in(reg_weight_3_23), .partial_sum_in(reg_psum_3_23), .reg_activation(reg_activation_4_23), .reg_weight(reg_weight_4_23), .reg_partial_sum(reg_psum_4_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_24( .activation_in(reg_activation_4_23), .weight_in(reg_weight_3_24), .partial_sum_in(reg_psum_3_24), .reg_activation(reg_activation_4_24), .reg_weight(reg_weight_4_24), .reg_partial_sum(reg_psum_4_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_25( .activation_in(reg_activation_4_24), .weight_in(reg_weight_3_25), .partial_sum_in(reg_psum_3_25), .reg_activation(reg_activation_4_25), .reg_weight(reg_weight_4_25), .reg_partial_sum(reg_psum_4_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_26( .activation_in(reg_activation_4_25), .weight_in(reg_weight_3_26), .partial_sum_in(reg_psum_3_26), .reg_activation(reg_activation_4_26), .reg_weight(reg_weight_4_26), .reg_partial_sum(reg_psum_4_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_27( .activation_in(reg_activation_4_26), .weight_in(reg_weight_3_27), .partial_sum_in(reg_psum_3_27), .reg_activation(reg_activation_4_27), .reg_weight(reg_weight_4_27), .reg_partial_sum(reg_psum_4_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_28( .activation_in(reg_activation_4_27), .weight_in(reg_weight_3_28), .partial_sum_in(reg_psum_3_28), .reg_activation(reg_activation_4_28), .reg_weight(reg_weight_4_28), .reg_partial_sum(reg_psum_4_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_29( .activation_in(reg_activation_4_28), .weight_in(reg_weight_3_29), .partial_sum_in(reg_psum_3_29), .reg_activation(reg_activation_4_29), .reg_weight(reg_weight_4_29), .reg_partial_sum(reg_psum_4_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_30( .activation_in(reg_activation_4_29), .weight_in(reg_weight_3_30), .partial_sum_in(reg_psum_3_30), .reg_activation(reg_activation_4_30), .reg_weight(reg_weight_4_30), .reg_partial_sum(reg_psum_4_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_31( .activation_in(reg_activation_4_30), .weight_in(reg_weight_3_31), .partial_sum_in(reg_psum_3_31), .reg_activation(reg_activation_4_31), .reg_weight(reg_weight_4_31), .reg_partial_sum(reg_psum_4_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_32( .activation_in(reg_activation_4_31), .weight_in(reg_weight_3_32), .partial_sum_in(reg_psum_3_32), .reg_activation(reg_activation_4_32), .reg_weight(reg_weight_4_32), .reg_partial_sum(reg_psum_4_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_33( .activation_in(reg_activation_4_32), .weight_in(reg_weight_3_33), .partial_sum_in(reg_psum_3_33), .reg_activation(reg_activation_4_33), .reg_weight(reg_weight_4_33), .reg_partial_sum(reg_psum_4_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_34( .activation_in(reg_activation_4_33), .weight_in(reg_weight_3_34), .partial_sum_in(reg_psum_3_34), .reg_activation(reg_activation_4_34), .reg_weight(reg_weight_4_34), .reg_partial_sum(reg_psum_4_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_35( .activation_in(reg_activation_4_34), .weight_in(reg_weight_3_35), .partial_sum_in(reg_psum_3_35), .reg_activation(reg_activation_4_35), .reg_weight(reg_weight_4_35), .reg_partial_sum(reg_psum_4_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_36( .activation_in(reg_activation_4_35), .weight_in(reg_weight_3_36), .partial_sum_in(reg_psum_3_36), .reg_activation(reg_activation_4_36), .reg_weight(reg_weight_4_36), .reg_partial_sum(reg_psum_4_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_37( .activation_in(reg_activation_4_36), .weight_in(reg_weight_3_37), .partial_sum_in(reg_psum_3_37), .reg_activation(reg_activation_4_37), .reg_weight(reg_weight_4_37), .reg_partial_sum(reg_psum_4_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_38( .activation_in(reg_activation_4_37), .weight_in(reg_weight_3_38), .partial_sum_in(reg_psum_3_38), .reg_activation(reg_activation_4_38), .reg_weight(reg_weight_4_38), .reg_partial_sum(reg_psum_4_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_39( .activation_in(reg_activation_4_38), .weight_in(reg_weight_3_39), .partial_sum_in(reg_psum_3_39), .reg_activation(reg_activation_4_39), .reg_weight(reg_weight_4_39), .reg_partial_sum(reg_psum_4_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_40( .activation_in(reg_activation_4_39), .weight_in(reg_weight_3_40), .partial_sum_in(reg_psum_3_40), .reg_activation(reg_activation_4_40), .reg_weight(reg_weight_4_40), .reg_partial_sum(reg_psum_4_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_41( .activation_in(reg_activation_4_40), .weight_in(reg_weight_3_41), .partial_sum_in(reg_psum_3_41), .reg_activation(reg_activation_4_41), .reg_weight(reg_weight_4_41), .reg_partial_sum(reg_psum_4_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_42( .activation_in(reg_activation_4_41), .weight_in(reg_weight_3_42), .partial_sum_in(reg_psum_3_42), .reg_activation(reg_activation_4_42), .reg_weight(reg_weight_4_42), .reg_partial_sum(reg_psum_4_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_43( .activation_in(reg_activation_4_42), .weight_in(reg_weight_3_43), .partial_sum_in(reg_psum_3_43), .reg_activation(reg_activation_4_43), .reg_weight(reg_weight_4_43), .reg_partial_sum(reg_psum_4_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_44( .activation_in(reg_activation_4_43), .weight_in(reg_weight_3_44), .partial_sum_in(reg_psum_3_44), .reg_activation(reg_activation_4_44), .reg_weight(reg_weight_4_44), .reg_partial_sum(reg_psum_4_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_45( .activation_in(reg_activation_4_44), .weight_in(reg_weight_3_45), .partial_sum_in(reg_psum_3_45), .reg_activation(reg_activation_4_45), .reg_weight(reg_weight_4_45), .reg_partial_sum(reg_psum_4_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_46( .activation_in(reg_activation_4_45), .weight_in(reg_weight_3_46), .partial_sum_in(reg_psum_3_46), .reg_activation(reg_activation_4_46), .reg_weight(reg_weight_4_46), .reg_partial_sum(reg_psum_4_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_47( .activation_in(reg_activation_4_46), .weight_in(reg_weight_3_47), .partial_sum_in(reg_psum_3_47), .reg_activation(reg_activation_4_47), .reg_weight(reg_weight_4_47), .reg_partial_sum(reg_psum_4_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_48( .activation_in(reg_activation_4_47), .weight_in(reg_weight_3_48), .partial_sum_in(reg_psum_3_48), .reg_activation(reg_activation_4_48), .reg_weight(reg_weight_4_48), .reg_partial_sum(reg_psum_4_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_49( .activation_in(reg_activation_4_48), .weight_in(reg_weight_3_49), .partial_sum_in(reg_psum_3_49), .reg_activation(reg_activation_4_49), .reg_weight(reg_weight_4_49), .reg_partial_sum(reg_psum_4_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_50( .activation_in(reg_activation_4_49), .weight_in(reg_weight_3_50), .partial_sum_in(reg_psum_3_50), .reg_activation(reg_activation_4_50), .reg_weight(reg_weight_4_50), .reg_partial_sum(reg_psum_4_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_51( .activation_in(reg_activation_4_50), .weight_in(reg_weight_3_51), .partial_sum_in(reg_psum_3_51), .reg_activation(reg_activation_4_51), .reg_weight(reg_weight_4_51), .reg_partial_sum(reg_psum_4_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_52( .activation_in(reg_activation_4_51), .weight_in(reg_weight_3_52), .partial_sum_in(reg_psum_3_52), .reg_activation(reg_activation_4_52), .reg_weight(reg_weight_4_52), .reg_partial_sum(reg_psum_4_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_53( .activation_in(reg_activation_4_52), .weight_in(reg_weight_3_53), .partial_sum_in(reg_psum_3_53), .reg_activation(reg_activation_4_53), .reg_weight(reg_weight_4_53), .reg_partial_sum(reg_psum_4_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_54( .activation_in(reg_activation_4_53), .weight_in(reg_weight_3_54), .partial_sum_in(reg_psum_3_54), .reg_activation(reg_activation_4_54), .reg_weight(reg_weight_4_54), .reg_partial_sum(reg_psum_4_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_55( .activation_in(reg_activation_4_54), .weight_in(reg_weight_3_55), .partial_sum_in(reg_psum_3_55), .reg_activation(reg_activation_4_55), .reg_weight(reg_weight_4_55), .reg_partial_sum(reg_psum_4_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_56( .activation_in(reg_activation_4_55), .weight_in(reg_weight_3_56), .partial_sum_in(reg_psum_3_56), .reg_activation(reg_activation_4_56), .reg_weight(reg_weight_4_56), .reg_partial_sum(reg_psum_4_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_57( .activation_in(reg_activation_4_56), .weight_in(reg_weight_3_57), .partial_sum_in(reg_psum_3_57), .reg_activation(reg_activation_4_57), .reg_weight(reg_weight_4_57), .reg_partial_sum(reg_psum_4_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_58( .activation_in(reg_activation_4_57), .weight_in(reg_weight_3_58), .partial_sum_in(reg_psum_3_58), .reg_activation(reg_activation_4_58), .reg_weight(reg_weight_4_58), .reg_partial_sum(reg_psum_4_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_59( .activation_in(reg_activation_4_58), .weight_in(reg_weight_3_59), .partial_sum_in(reg_psum_3_59), .reg_activation(reg_activation_4_59), .reg_weight(reg_weight_4_59), .reg_partial_sum(reg_psum_4_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_60( .activation_in(reg_activation_4_59), .weight_in(reg_weight_3_60), .partial_sum_in(reg_psum_3_60), .reg_activation(reg_activation_4_60), .reg_weight(reg_weight_4_60), .reg_partial_sum(reg_psum_4_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_61( .activation_in(reg_activation_4_60), .weight_in(reg_weight_3_61), .partial_sum_in(reg_psum_3_61), .reg_activation(reg_activation_4_61), .reg_weight(reg_weight_4_61), .reg_partial_sum(reg_psum_4_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_62( .activation_in(reg_activation_4_61), .weight_in(reg_weight_3_62), .partial_sum_in(reg_psum_3_62), .reg_activation(reg_activation_4_62), .reg_weight(reg_weight_4_62), .reg_partial_sum(reg_psum_4_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_63( .activation_in(reg_activation_4_62), .weight_in(reg_weight_3_63), .partial_sum_in(reg_psum_3_63), .reg_weight(reg_weight_4_63), .reg_partial_sum(reg_psum_4_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_0( .activation_in(in_activation_5), .weight_in(reg_weight_4_0), .partial_sum_in(reg_psum_4_0), .reg_activation(reg_activation_5_0), .reg_weight(reg_weight_5_0), .reg_partial_sum(reg_psum_5_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_1( .activation_in(reg_activation_5_0), .weight_in(reg_weight_4_1), .partial_sum_in(reg_psum_4_1), .reg_activation(reg_activation_5_1), .reg_weight(reg_weight_5_1), .reg_partial_sum(reg_psum_5_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_2( .activation_in(reg_activation_5_1), .weight_in(reg_weight_4_2), .partial_sum_in(reg_psum_4_2), .reg_activation(reg_activation_5_2), .reg_weight(reg_weight_5_2), .reg_partial_sum(reg_psum_5_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_3( .activation_in(reg_activation_5_2), .weight_in(reg_weight_4_3), .partial_sum_in(reg_psum_4_3), .reg_activation(reg_activation_5_3), .reg_weight(reg_weight_5_3), .reg_partial_sum(reg_psum_5_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_4( .activation_in(reg_activation_5_3), .weight_in(reg_weight_4_4), .partial_sum_in(reg_psum_4_4), .reg_activation(reg_activation_5_4), .reg_weight(reg_weight_5_4), .reg_partial_sum(reg_psum_5_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_5( .activation_in(reg_activation_5_4), .weight_in(reg_weight_4_5), .partial_sum_in(reg_psum_4_5), .reg_activation(reg_activation_5_5), .reg_weight(reg_weight_5_5), .reg_partial_sum(reg_psum_5_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_6( .activation_in(reg_activation_5_5), .weight_in(reg_weight_4_6), .partial_sum_in(reg_psum_4_6), .reg_activation(reg_activation_5_6), .reg_weight(reg_weight_5_6), .reg_partial_sum(reg_psum_5_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_7( .activation_in(reg_activation_5_6), .weight_in(reg_weight_4_7), .partial_sum_in(reg_psum_4_7), .reg_activation(reg_activation_5_7), .reg_weight(reg_weight_5_7), .reg_partial_sum(reg_psum_5_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_8( .activation_in(reg_activation_5_7), .weight_in(reg_weight_4_8), .partial_sum_in(reg_psum_4_8), .reg_activation(reg_activation_5_8), .reg_weight(reg_weight_5_8), .reg_partial_sum(reg_psum_5_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_9( .activation_in(reg_activation_5_8), .weight_in(reg_weight_4_9), .partial_sum_in(reg_psum_4_9), .reg_activation(reg_activation_5_9), .reg_weight(reg_weight_5_9), .reg_partial_sum(reg_psum_5_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_10( .activation_in(reg_activation_5_9), .weight_in(reg_weight_4_10), .partial_sum_in(reg_psum_4_10), .reg_activation(reg_activation_5_10), .reg_weight(reg_weight_5_10), .reg_partial_sum(reg_psum_5_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_11( .activation_in(reg_activation_5_10), .weight_in(reg_weight_4_11), .partial_sum_in(reg_psum_4_11), .reg_activation(reg_activation_5_11), .reg_weight(reg_weight_5_11), .reg_partial_sum(reg_psum_5_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_12( .activation_in(reg_activation_5_11), .weight_in(reg_weight_4_12), .partial_sum_in(reg_psum_4_12), .reg_activation(reg_activation_5_12), .reg_weight(reg_weight_5_12), .reg_partial_sum(reg_psum_5_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_13( .activation_in(reg_activation_5_12), .weight_in(reg_weight_4_13), .partial_sum_in(reg_psum_4_13), .reg_activation(reg_activation_5_13), .reg_weight(reg_weight_5_13), .reg_partial_sum(reg_psum_5_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_14( .activation_in(reg_activation_5_13), .weight_in(reg_weight_4_14), .partial_sum_in(reg_psum_4_14), .reg_activation(reg_activation_5_14), .reg_weight(reg_weight_5_14), .reg_partial_sum(reg_psum_5_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_15( .activation_in(reg_activation_5_14), .weight_in(reg_weight_4_15), .partial_sum_in(reg_psum_4_15), .reg_activation(reg_activation_5_15), .reg_weight(reg_weight_5_15), .reg_partial_sum(reg_psum_5_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_16( .activation_in(reg_activation_5_15), .weight_in(reg_weight_4_16), .partial_sum_in(reg_psum_4_16), .reg_activation(reg_activation_5_16), .reg_weight(reg_weight_5_16), .reg_partial_sum(reg_psum_5_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_17( .activation_in(reg_activation_5_16), .weight_in(reg_weight_4_17), .partial_sum_in(reg_psum_4_17), .reg_activation(reg_activation_5_17), .reg_weight(reg_weight_5_17), .reg_partial_sum(reg_psum_5_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_18( .activation_in(reg_activation_5_17), .weight_in(reg_weight_4_18), .partial_sum_in(reg_psum_4_18), .reg_activation(reg_activation_5_18), .reg_weight(reg_weight_5_18), .reg_partial_sum(reg_psum_5_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_19( .activation_in(reg_activation_5_18), .weight_in(reg_weight_4_19), .partial_sum_in(reg_psum_4_19), .reg_activation(reg_activation_5_19), .reg_weight(reg_weight_5_19), .reg_partial_sum(reg_psum_5_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_20( .activation_in(reg_activation_5_19), .weight_in(reg_weight_4_20), .partial_sum_in(reg_psum_4_20), .reg_activation(reg_activation_5_20), .reg_weight(reg_weight_5_20), .reg_partial_sum(reg_psum_5_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_21( .activation_in(reg_activation_5_20), .weight_in(reg_weight_4_21), .partial_sum_in(reg_psum_4_21), .reg_activation(reg_activation_5_21), .reg_weight(reg_weight_5_21), .reg_partial_sum(reg_psum_5_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_22( .activation_in(reg_activation_5_21), .weight_in(reg_weight_4_22), .partial_sum_in(reg_psum_4_22), .reg_activation(reg_activation_5_22), .reg_weight(reg_weight_5_22), .reg_partial_sum(reg_psum_5_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_23( .activation_in(reg_activation_5_22), .weight_in(reg_weight_4_23), .partial_sum_in(reg_psum_4_23), .reg_activation(reg_activation_5_23), .reg_weight(reg_weight_5_23), .reg_partial_sum(reg_psum_5_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_24( .activation_in(reg_activation_5_23), .weight_in(reg_weight_4_24), .partial_sum_in(reg_psum_4_24), .reg_activation(reg_activation_5_24), .reg_weight(reg_weight_5_24), .reg_partial_sum(reg_psum_5_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_25( .activation_in(reg_activation_5_24), .weight_in(reg_weight_4_25), .partial_sum_in(reg_psum_4_25), .reg_activation(reg_activation_5_25), .reg_weight(reg_weight_5_25), .reg_partial_sum(reg_psum_5_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_26( .activation_in(reg_activation_5_25), .weight_in(reg_weight_4_26), .partial_sum_in(reg_psum_4_26), .reg_activation(reg_activation_5_26), .reg_weight(reg_weight_5_26), .reg_partial_sum(reg_psum_5_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_27( .activation_in(reg_activation_5_26), .weight_in(reg_weight_4_27), .partial_sum_in(reg_psum_4_27), .reg_activation(reg_activation_5_27), .reg_weight(reg_weight_5_27), .reg_partial_sum(reg_psum_5_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_28( .activation_in(reg_activation_5_27), .weight_in(reg_weight_4_28), .partial_sum_in(reg_psum_4_28), .reg_activation(reg_activation_5_28), .reg_weight(reg_weight_5_28), .reg_partial_sum(reg_psum_5_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_29( .activation_in(reg_activation_5_28), .weight_in(reg_weight_4_29), .partial_sum_in(reg_psum_4_29), .reg_activation(reg_activation_5_29), .reg_weight(reg_weight_5_29), .reg_partial_sum(reg_psum_5_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_30( .activation_in(reg_activation_5_29), .weight_in(reg_weight_4_30), .partial_sum_in(reg_psum_4_30), .reg_activation(reg_activation_5_30), .reg_weight(reg_weight_5_30), .reg_partial_sum(reg_psum_5_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_31( .activation_in(reg_activation_5_30), .weight_in(reg_weight_4_31), .partial_sum_in(reg_psum_4_31), .reg_activation(reg_activation_5_31), .reg_weight(reg_weight_5_31), .reg_partial_sum(reg_psum_5_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_32( .activation_in(reg_activation_5_31), .weight_in(reg_weight_4_32), .partial_sum_in(reg_psum_4_32), .reg_activation(reg_activation_5_32), .reg_weight(reg_weight_5_32), .reg_partial_sum(reg_psum_5_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_33( .activation_in(reg_activation_5_32), .weight_in(reg_weight_4_33), .partial_sum_in(reg_psum_4_33), .reg_activation(reg_activation_5_33), .reg_weight(reg_weight_5_33), .reg_partial_sum(reg_psum_5_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_34( .activation_in(reg_activation_5_33), .weight_in(reg_weight_4_34), .partial_sum_in(reg_psum_4_34), .reg_activation(reg_activation_5_34), .reg_weight(reg_weight_5_34), .reg_partial_sum(reg_psum_5_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_35( .activation_in(reg_activation_5_34), .weight_in(reg_weight_4_35), .partial_sum_in(reg_psum_4_35), .reg_activation(reg_activation_5_35), .reg_weight(reg_weight_5_35), .reg_partial_sum(reg_psum_5_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_36( .activation_in(reg_activation_5_35), .weight_in(reg_weight_4_36), .partial_sum_in(reg_psum_4_36), .reg_activation(reg_activation_5_36), .reg_weight(reg_weight_5_36), .reg_partial_sum(reg_psum_5_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_37( .activation_in(reg_activation_5_36), .weight_in(reg_weight_4_37), .partial_sum_in(reg_psum_4_37), .reg_activation(reg_activation_5_37), .reg_weight(reg_weight_5_37), .reg_partial_sum(reg_psum_5_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_38( .activation_in(reg_activation_5_37), .weight_in(reg_weight_4_38), .partial_sum_in(reg_psum_4_38), .reg_activation(reg_activation_5_38), .reg_weight(reg_weight_5_38), .reg_partial_sum(reg_psum_5_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_39( .activation_in(reg_activation_5_38), .weight_in(reg_weight_4_39), .partial_sum_in(reg_psum_4_39), .reg_activation(reg_activation_5_39), .reg_weight(reg_weight_5_39), .reg_partial_sum(reg_psum_5_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_40( .activation_in(reg_activation_5_39), .weight_in(reg_weight_4_40), .partial_sum_in(reg_psum_4_40), .reg_activation(reg_activation_5_40), .reg_weight(reg_weight_5_40), .reg_partial_sum(reg_psum_5_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_41( .activation_in(reg_activation_5_40), .weight_in(reg_weight_4_41), .partial_sum_in(reg_psum_4_41), .reg_activation(reg_activation_5_41), .reg_weight(reg_weight_5_41), .reg_partial_sum(reg_psum_5_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_42( .activation_in(reg_activation_5_41), .weight_in(reg_weight_4_42), .partial_sum_in(reg_psum_4_42), .reg_activation(reg_activation_5_42), .reg_weight(reg_weight_5_42), .reg_partial_sum(reg_psum_5_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_43( .activation_in(reg_activation_5_42), .weight_in(reg_weight_4_43), .partial_sum_in(reg_psum_4_43), .reg_activation(reg_activation_5_43), .reg_weight(reg_weight_5_43), .reg_partial_sum(reg_psum_5_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_44( .activation_in(reg_activation_5_43), .weight_in(reg_weight_4_44), .partial_sum_in(reg_psum_4_44), .reg_activation(reg_activation_5_44), .reg_weight(reg_weight_5_44), .reg_partial_sum(reg_psum_5_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_45( .activation_in(reg_activation_5_44), .weight_in(reg_weight_4_45), .partial_sum_in(reg_psum_4_45), .reg_activation(reg_activation_5_45), .reg_weight(reg_weight_5_45), .reg_partial_sum(reg_psum_5_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_46( .activation_in(reg_activation_5_45), .weight_in(reg_weight_4_46), .partial_sum_in(reg_psum_4_46), .reg_activation(reg_activation_5_46), .reg_weight(reg_weight_5_46), .reg_partial_sum(reg_psum_5_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_47( .activation_in(reg_activation_5_46), .weight_in(reg_weight_4_47), .partial_sum_in(reg_psum_4_47), .reg_activation(reg_activation_5_47), .reg_weight(reg_weight_5_47), .reg_partial_sum(reg_psum_5_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_48( .activation_in(reg_activation_5_47), .weight_in(reg_weight_4_48), .partial_sum_in(reg_psum_4_48), .reg_activation(reg_activation_5_48), .reg_weight(reg_weight_5_48), .reg_partial_sum(reg_psum_5_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_49( .activation_in(reg_activation_5_48), .weight_in(reg_weight_4_49), .partial_sum_in(reg_psum_4_49), .reg_activation(reg_activation_5_49), .reg_weight(reg_weight_5_49), .reg_partial_sum(reg_psum_5_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_50( .activation_in(reg_activation_5_49), .weight_in(reg_weight_4_50), .partial_sum_in(reg_psum_4_50), .reg_activation(reg_activation_5_50), .reg_weight(reg_weight_5_50), .reg_partial_sum(reg_psum_5_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_51( .activation_in(reg_activation_5_50), .weight_in(reg_weight_4_51), .partial_sum_in(reg_psum_4_51), .reg_activation(reg_activation_5_51), .reg_weight(reg_weight_5_51), .reg_partial_sum(reg_psum_5_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_52( .activation_in(reg_activation_5_51), .weight_in(reg_weight_4_52), .partial_sum_in(reg_psum_4_52), .reg_activation(reg_activation_5_52), .reg_weight(reg_weight_5_52), .reg_partial_sum(reg_psum_5_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_53( .activation_in(reg_activation_5_52), .weight_in(reg_weight_4_53), .partial_sum_in(reg_psum_4_53), .reg_activation(reg_activation_5_53), .reg_weight(reg_weight_5_53), .reg_partial_sum(reg_psum_5_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_54( .activation_in(reg_activation_5_53), .weight_in(reg_weight_4_54), .partial_sum_in(reg_psum_4_54), .reg_activation(reg_activation_5_54), .reg_weight(reg_weight_5_54), .reg_partial_sum(reg_psum_5_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_55( .activation_in(reg_activation_5_54), .weight_in(reg_weight_4_55), .partial_sum_in(reg_psum_4_55), .reg_activation(reg_activation_5_55), .reg_weight(reg_weight_5_55), .reg_partial_sum(reg_psum_5_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_56( .activation_in(reg_activation_5_55), .weight_in(reg_weight_4_56), .partial_sum_in(reg_psum_4_56), .reg_activation(reg_activation_5_56), .reg_weight(reg_weight_5_56), .reg_partial_sum(reg_psum_5_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_57( .activation_in(reg_activation_5_56), .weight_in(reg_weight_4_57), .partial_sum_in(reg_psum_4_57), .reg_activation(reg_activation_5_57), .reg_weight(reg_weight_5_57), .reg_partial_sum(reg_psum_5_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_58( .activation_in(reg_activation_5_57), .weight_in(reg_weight_4_58), .partial_sum_in(reg_psum_4_58), .reg_activation(reg_activation_5_58), .reg_weight(reg_weight_5_58), .reg_partial_sum(reg_psum_5_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_59( .activation_in(reg_activation_5_58), .weight_in(reg_weight_4_59), .partial_sum_in(reg_psum_4_59), .reg_activation(reg_activation_5_59), .reg_weight(reg_weight_5_59), .reg_partial_sum(reg_psum_5_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_60( .activation_in(reg_activation_5_59), .weight_in(reg_weight_4_60), .partial_sum_in(reg_psum_4_60), .reg_activation(reg_activation_5_60), .reg_weight(reg_weight_5_60), .reg_partial_sum(reg_psum_5_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_61( .activation_in(reg_activation_5_60), .weight_in(reg_weight_4_61), .partial_sum_in(reg_psum_4_61), .reg_activation(reg_activation_5_61), .reg_weight(reg_weight_5_61), .reg_partial_sum(reg_psum_5_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_62( .activation_in(reg_activation_5_61), .weight_in(reg_weight_4_62), .partial_sum_in(reg_psum_4_62), .reg_activation(reg_activation_5_62), .reg_weight(reg_weight_5_62), .reg_partial_sum(reg_psum_5_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_63( .activation_in(reg_activation_5_62), .weight_in(reg_weight_4_63), .partial_sum_in(reg_psum_4_63), .reg_weight(reg_weight_5_63), .reg_partial_sum(reg_psum_5_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_0( .activation_in(in_activation_6), .weight_in(reg_weight_5_0), .partial_sum_in(reg_psum_5_0), .reg_activation(reg_activation_6_0), .reg_weight(reg_weight_6_0), .reg_partial_sum(reg_psum_6_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_1( .activation_in(reg_activation_6_0), .weight_in(reg_weight_5_1), .partial_sum_in(reg_psum_5_1), .reg_activation(reg_activation_6_1), .reg_weight(reg_weight_6_1), .reg_partial_sum(reg_psum_6_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_2( .activation_in(reg_activation_6_1), .weight_in(reg_weight_5_2), .partial_sum_in(reg_psum_5_2), .reg_activation(reg_activation_6_2), .reg_weight(reg_weight_6_2), .reg_partial_sum(reg_psum_6_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_3( .activation_in(reg_activation_6_2), .weight_in(reg_weight_5_3), .partial_sum_in(reg_psum_5_3), .reg_activation(reg_activation_6_3), .reg_weight(reg_weight_6_3), .reg_partial_sum(reg_psum_6_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_4( .activation_in(reg_activation_6_3), .weight_in(reg_weight_5_4), .partial_sum_in(reg_psum_5_4), .reg_activation(reg_activation_6_4), .reg_weight(reg_weight_6_4), .reg_partial_sum(reg_psum_6_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_5( .activation_in(reg_activation_6_4), .weight_in(reg_weight_5_5), .partial_sum_in(reg_psum_5_5), .reg_activation(reg_activation_6_5), .reg_weight(reg_weight_6_5), .reg_partial_sum(reg_psum_6_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_6( .activation_in(reg_activation_6_5), .weight_in(reg_weight_5_6), .partial_sum_in(reg_psum_5_6), .reg_activation(reg_activation_6_6), .reg_weight(reg_weight_6_6), .reg_partial_sum(reg_psum_6_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_7( .activation_in(reg_activation_6_6), .weight_in(reg_weight_5_7), .partial_sum_in(reg_psum_5_7), .reg_activation(reg_activation_6_7), .reg_weight(reg_weight_6_7), .reg_partial_sum(reg_psum_6_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_8( .activation_in(reg_activation_6_7), .weight_in(reg_weight_5_8), .partial_sum_in(reg_psum_5_8), .reg_activation(reg_activation_6_8), .reg_weight(reg_weight_6_8), .reg_partial_sum(reg_psum_6_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_9( .activation_in(reg_activation_6_8), .weight_in(reg_weight_5_9), .partial_sum_in(reg_psum_5_9), .reg_activation(reg_activation_6_9), .reg_weight(reg_weight_6_9), .reg_partial_sum(reg_psum_6_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_10( .activation_in(reg_activation_6_9), .weight_in(reg_weight_5_10), .partial_sum_in(reg_psum_5_10), .reg_activation(reg_activation_6_10), .reg_weight(reg_weight_6_10), .reg_partial_sum(reg_psum_6_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_11( .activation_in(reg_activation_6_10), .weight_in(reg_weight_5_11), .partial_sum_in(reg_psum_5_11), .reg_activation(reg_activation_6_11), .reg_weight(reg_weight_6_11), .reg_partial_sum(reg_psum_6_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_12( .activation_in(reg_activation_6_11), .weight_in(reg_weight_5_12), .partial_sum_in(reg_psum_5_12), .reg_activation(reg_activation_6_12), .reg_weight(reg_weight_6_12), .reg_partial_sum(reg_psum_6_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_13( .activation_in(reg_activation_6_12), .weight_in(reg_weight_5_13), .partial_sum_in(reg_psum_5_13), .reg_activation(reg_activation_6_13), .reg_weight(reg_weight_6_13), .reg_partial_sum(reg_psum_6_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_14( .activation_in(reg_activation_6_13), .weight_in(reg_weight_5_14), .partial_sum_in(reg_psum_5_14), .reg_activation(reg_activation_6_14), .reg_weight(reg_weight_6_14), .reg_partial_sum(reg_psum_6_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_15( .activation_in(reg_activation_6_14), .weight_in(reg_weight_5_15), .partial_sum_in(reg_psum_5_15), .reg_activation(reg_activation_6_15), .reg_weight(reg_weight_6_15), .reg_partial_sum(reg_psum_6_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_16( .activation_in(reg_activation_6_15), .weight_in(reg_weight_5_16), .partial_sum_in(reg_psum_5_16), .reg_activation(reg_activation_6_16), .reg_weight(reg_weight_6_16), .reg_partial_sum(reg_psum_6_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_17( .activation_in(reg_activation_6_16), .weight_in(reg_weight_5_17), .partial_sum_in(reg_psum_5_17), .reg_activation(reg_activation_6_17), .reg_weight(reg_weight_6_17), .reg_partial_sum(reg_psum_6_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_18( .activation_in(reg_activation_6_17), .weight_in(reg_weight_5_18), .partial_sum_in(reg_psum_5_18), .reg_activation(reg_activation_6_18), .reg_weight(reg_weight_6_18), .reg_partial_sum(reg_psum_6_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_19( .activation_in(reg_activation_6_18), .weight_in(reg_weight_5_19), .partial_sum_in(reg_psum_5_19), .reg_activation(reg_activation_6_19), .reg_weight(reg_weight_6_19), .reg_partial_sum(reg_psum_6_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_20( .activation_in(reg_activation_6_19), .weight_in(reg_weight_5_20), .partial_sum_in(reg_psum_5_20), .reg_activation(reg_activation_6_20), .reg_weight(reg_weight_6_20), .reg_partial_sum(reg_psum_6_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_21( .activation_in(reg_activation_6_20), .weight_in(reg_weight_5_21), .partial_sum_in(reg_psum_5_21), .reg_activation(reg_activation_6_21), .reg_weight(reg_weight_6_21), .reg_partial_sum(reg_psum_6_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_22( .activation_in(reg_activation_6_21), .weight_in(reg_weight_5_22), .partial_sum_in(reg_psum_5_22), .reg_activation(reg_activation_6_22), .reg_weight(reg_weight_6_22), .reg_partial_sum(reg_psum_6_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_23( .activation_in(reg_activation_6_22), .weight_in(reg_weight_5_23), .partial_sum_in(reg_psum_5_23), .reg_activation(reg_activation_6_23), .reg_weight(reg_weight_6_23), .reg_partial_sum(reg_psum_6_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_24( .activation_in(reg_activation_6_23), .weight_in(reg_weight_5_24), .partial_sum_in(reg_psum_5_24), .reg_activation(reg_activation_6_24), .reg_weight(reg_weight_6_24), .reg_partial_sum(reg_psum_6_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_25( .activation_in(reg_activation_6_24), .weight_in(reg_weight_5_25), .partial_sum_in(reg_psum_5_25), .reg_activation(reg_activation_6_25), .reg_weight(reg_weight_6_25), .reg_partial_sum(reg_psum_6_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_26( .activation_in(reg_activation_6_25), .weight_in(reg_weight_5_26), .partial_sum_in(reg_psum_5_26), .reg_activation(reg_activation_6_26), .reg_weight(reg_weight_6_26), .reg_partial_sum(reg_psum_6_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_27( .activation_in(reg_activation_6_26), .weight_in(reg_weight_5_27), .partial_sum_in(reg_psum_5_27), .reg_activation(reg_activation_6_27), .reg_weight(reg_weight_6_27), .reg_partial_sum(reg_psum_6_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_28( .activation_in(reg_activation_6_27), .weight_in(reg_weight_5_28), .partial_sum_in(reg_psum_5_28), .reg_activation(reg_activation_6_28), .reg_weight(reg_weight_6_28), .reg_partial_sum(reg_psum_6_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_29( .activation_in(reg_activation_6_28), .weight_in(reg_weight_5_29), .partial_sum_in(reg_psum_5_29), .reg_activation(reg_activation_6_29), .reg_weight(reg_weight_6_29), .reg_partial_sum(reg_psum_6_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_30( .activation_in(reg_activation_6_29), .weight_in(reg_weight_5_30), .partial_sum_in(reg_psum_5_30), .reg_activation(reg_activation_6_30), .reg_weight(reg_weight_6_30), .reg_partial_sum(reg_psum_6_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_31( .activation_in(reg_activation_6_30), .weight_in(reg_weight_5_31), .partial_sum_in(reg_psum_5_31), .reg_activation(reg_activation_6_31), .reg_weight(reg_weight_6_31), .reg_partial_sum(reg_psum_6_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_32( .activation_in(reg_activation_6_31), .weight_in(reg_weight_5_32), .partial_sum_in(reg_psum_5_32), .reg_activation(reg_activation_6_32), .reg_weight(reg_weight_6_32), .reg_partial_sum(reg_psum_6_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_33( .activation_in(reg_activation_6_32), .weight_in(reg_weight_5_33), .partial_sum_in(reg_psum_5_33), .reg_activation(reg_activation_6_33), .reg_weight(reg_weight_6_33), .reg_partial_sum(reg_psum_6_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_34( .activation_in(reg_activation_6_33), .weight_in(reg_weight_5_34), .partial_sum_in(reg_psum_5_34), .reg_activation(reg_activation_6_34), .reg_weight(reg_weight_6_34), .reg_partial_sum(reg_psum_6_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_35( .activation_in(reg_activation_6_34), .weight_in(reg_weight_5_35), .partial_sum_in(reg_psum_5_35), .reg_activation(reg_activation_6_35), .reg_weight(reg_weight_6_35), .reg_partial_sum(reg_psum_6_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_36( .activation_in(reg_activation_6_35), .weight_in(reg_weight_5_36), .partial_sum_in(reg_psum_5_36), .reg_activation(reg_activation_6_36), .reg_weight(reg_weight_6_36), .reg_partial_sum(reg_psum_6_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_37( .activation_in(reg_activation_6_36), .weight_in(reg_weight_5_37), .partial_sum_in(reg_psum_5_37), .reg_activation(reg_activation_6_37), .reg_weight(reg_weight_6_37), .reg_partial_sum(reg_psum_6_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_38( .activation_in(reg_activation_6_37), .weight_in(reg_weight_5_38), .partial_sum_in(reg_psum_5_38), .reg_activation(reg_activation_6_38), .reg_weight(reg_weight_6_38), .reg_partial_sum(reg_psum_6_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_39( .activation_in(reg_activation_6_38), .weight_in(reg_weight_5_39), .partial_sum_in(reg_psum_5_39), .reg_activation(reg_activation_6_39), .reg_weight(reg_weight_6_39), .reg_partial_sum(reg_psum_6_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_40( .activation_in(reg_activation_6_39), .weight_in(reg_weight_5_40), .partial_sum_in(reg_psum_5_40), .reg_activation(reg_activation_6_40), .reg_weight(reg_weight_6_40), .reg_partial_sum(reg_psum_6_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_41( .activation_in(reg_activation_6_40), .weight_in(reg_weight_5_41), .partial_sum_in(reg_psum_5_41), .reg_activation(reg_activation_6_41), .reg_weight(reg_weight_6_41), .reg_partial_sum(reg_psum_6_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_42( .activation_in(reg_activation_6_41), .weight_in(reg_weight_5_42), .partial_sum_in(reg_psum_5_42), .reg_activation(reg_activation_6_42), .reg_weight(reg_weight_6_42), .reg_partial_sum(reg_psum_6_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_43( .activation_in(reg_activation_6_42), .weight_in(reg_weight_5_43), .partial_sum_in(reg_psum_5_43), .reg_activation(reg_activation_6_43), .reg_weight(reg_weight_6_43), .reg_partial_sum(reg_psum_6_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_44( .activation_in(reg_activation_6_43), .weight_in(reg_weight_5_44), .partial_sum_in(reg_psum_5_44), .reg_activation(reg_activation_6_44), .reg_weight(reg_weight_6_44), .reg_partial_sum(reg_psum_6_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_45( .activation_in(reg_activation_6_44), .weight_in(reg_weight_5_45), .partial_sum_in(reg_psum_5_45), .reg_activation(reg_activation_6_45), .reg_weight(reg_weight_6_45), .reg_partial_sum(reg_psum_6_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_46( .activation_in(reg_activation_6_45), .weight_in(reg_weight_5_46), .partial_sum_in(reg_psum_5_46), .reg_activation(reg_activation_6_46), .reg_weight(reg_weight_6_46), .reg_partial_sum(reg_psum_6_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_47( .activation_in(reg_activation_6_46), .weight_in(reg_weight_5_47), .partial_sum_in(reg_psum_5_47), .reg_activation(reg_activation_6_47), .reg_weight(reg_weight_6_47), .reg_partial_sum(reg_psum_6_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_48( .activation_in(reg_activation_6_47), .weight_in(reg_weight_5_48), .partial_sum_in(reg_psum_5_48), .reg_activation(reg_activation_6_48), .reg_weight(reg_weight_6_48), .reg_partial_sum(reg_psum_6_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_49( .activation_in(reg_activation_6_48), .weight_in(reg_weight_5_49), .partial_sum_in(reg_psum_5_49), .reg_activation(reg_activation_6_49), .reg_weight(reg_weight_6_49), .reg_partial_sum(reg_psum_6_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_50( .activation_in(reg_activation_6_49), .weight_in(reg_weight_5_50), .partial_sum_in(reg_psum_5_50), .reg_activation(reg_activation_6_50), .reg_weight(reg_weight_6_50), .reg_partial_sum(reg_psum_6_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_51( .activation_in(reg_activation_6_50), .weight_in(reg_weight_5_51), .partial_sum_in(reg_psum_5_51), .reg_activation(reg_activation_6_51), .reg_weight(reg_weight_6_51), .reg_partial_sum(reg_psum_6_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_52( .activation_in(reg_activation_6_51), .weight_in(reg_weight_5_52), .partial_sum_in(reg_psum_5_52), .reg_activation(reg_activation_6_52), .reg_weight(reg_weight_6_52), .reg_partial_sum(reg_psum_6_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_53( .activation_in(reg_activation_6_52), .weight_in(reg_weight_5_53), .partial_sum_in(reg_psum_5_53), .reg_activation(reg_activation_6_53), .reg_weight(reg_weight_6_53), .reg_partial_sum(reg_psum_6_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_54( .activation_in(reg_activation_6_53), .weight_in(reg_weight_5_54), .partial_sum_in(reg_psum_5_54), .reg_activation(reg_activation_6_54), .reg_weight(reg_weight_6_54), .reg_partial_sum(reg_psum_6_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_55( .activation_in(reg_activation_6_54), .weight_in(reg_weight_5_55), .partial_sum_in(reg_psum_5_55), .reg_activation(reg_activation_6_55), .reg_weight(reg_weight_6_55), .reg_partial_sum(reg_psum_6_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_56( .activation_in(reg_activation_6_55), .weight_in(reg_weight_5_56), .partial_sum_in(reg_psum_5_56), .reg_activation(reg_activation_6_56), .reg_weight(reg_weight_6_56), .reg_partial_sum(reg_psum_6_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_57( .activation_in(reg_activation_6_56), .weight_in(reg_weight_5_57), .partial_sum_in(reg_psum_5_57), .reg_activation(reg_activation_6_57), .reg_weight(reg_weight_6_57), .reg_partial_sum(reg_psum_6_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_58( .activation_in(reg_activation_6_57), .weight_in(reg_weight_5_58), .partial_sum_in(reg_psum_5_58), .reg_activation(reg_activation_6_58), .reg_weight(reg_weight_6_58), .reg_partial_sum(reg_psum_6_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_59( .activation_in(reg_activation_6_58), .weight_in(reg_weight_5_59), .partial_sum_in(reg_psum_5_59), .reg_activation(reg_activation_6_59), .reg_weight(reg_weight_6_59), .reg_partial_sum(reg_psum_6_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_60( .activation_in(reg_activation_6_59), .weight_in(reg_weight_5_60), .partial_sum_in(reg_psum_5_60), .reg_activation(reg_activation_6_60), .reg_weight(reg_weight_6_60), .reg_partial_sum(reg_psum_6_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_61( .activation_in(reg_activation_6_60), .weight_in(reg_weight_5_61), .partial_sum_in(reg_psum_5_61), .reg_activation(reg_activation_6_61), .reg_weight(reg_weight_6_61), .reg_partial_sum(reg_psum_6_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_62( .activation_in(reg_activation_6_61), .weight_in(reg_weight_5_62), .partial_sum_in(reg_psum_5_62), .reg_activation(reg_activation_6_62), .reg_weight(reg_weight_6_62), .reg_partial_sum(reg_psum_6_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_63( .activation_in(reg_activation_6_62), .weight_in(reg_weight_5_63), .partial_sum_in(reg_psum_5_63), .reg_weight(reg_weight_6_63), .reg_partial_sum(reg_psum_6_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_0( .activation_in(in_activation_7), .weight_in(reg_weight_6_0), .partial_sum_in(reg_psum_6_0), .reg_activation(reg_activation_7_0), .reg_weight(reg_weight_7_0), .reg_partial_sum(reg_psum_7_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_1( .activation_in(reg_activation_7_0), .weight_in(reg_weight_6_1), .partial_sum_in(reg_psum_6_1), .reg_activation(reg_activation_7_1), .reg_weight(reg_weight_7_1), .reg_partial_sum(reg_psum_7_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_2( .activation_in(reg_activation_7_1), .weight_in(reg_weight_6_2), .partial_sum_in(reg_psum_6_2), .reg_activation(reg_activation_7_2), .reg_weight(reg_weight_7_2), .reg_partial_sum(reg_psum_7_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_3( .activation_in(reg_activation_7_2), .weight_in(reg_weight_6_3), .partial_sum_in(reg_psum_6_3), .reg_activation(reg_activation_7_3), .reg_weight(reg_weight_7_3), .reg_partial_sum(reg_psum_7_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_4( .activation_in(reg_activation_7_3), .weight_in(reg_weight_6_4), .partial_sum_in(reg_psum_6_4), .reg_activation(reg_activation_7_4), .reg_weight(reg_weight_7_4), .reg_partial_sum(reg_psum_7_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_5( .activation_in(reg_activation_7_4), .weight_in(reg_weight_6_5), .partial_sum_in(reg_psum_6_5), .reg_activation(reg_activation_7_5), .reg_weight(reg_weight_7_5), .reg_partial_sum(reg_psum_7_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_6( .activation_in(reg_activation_7_5), .weight_in(reg_weight_6_6), .partial_sum_in(reg_psum_6_6), .reg_activation(reg_activation_7_6), .reg_weight(reg_weight_7_6), .reg_partial_sum(reg_psum_7_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_7( .activation_in(reg_activation_7_6), .weight_in(reg_weight_6_7), .partial_sum_in(reg_psum_6_7), .reg_activation(reg_activation_7_7), .reg_weight(reg_weight_7_7), .reg_partial_sum(reg_psum_7_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_8( .activation_in(reg_activation_7_7), .weight_in(reg_weight_6_8), .partial_sum_in(reg_psum_6_8), .reg_activation(reg_activation_7_8), .reg_weight(reg_weight_7_8), .reg_partial_sum(reg_psum_7_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_9( .activation_in(reg_activation_7_8), .weight_in(reg_weight_6_9), .partial_sum_in(reg_psum_6_9), .reg_activation(reg_activation_7_9), .reg_weight(reg_weight_7_9), .reg_partial_sum(reg_psum_7_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_10( .activation_in(reg_activation_7_9), .weight_in(reg_weight_6_10), .partial_sum_in(reg_psum_6_10), .reg_activation(reg_activation_7_10), .reg_weight(reg_weight_7_10), .reg_partial_sum(reg_psum_7_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_11( .activation_in(reg_activation_7_10), .weight_in(reg_weight_6_11), .partial_sum_in(reg_psum_6_11), .reg_activation(reg_activation_7_11), .reg_weight(reg_weight_7_11), .reg_partial_sum(reg_psum_7_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_12( .activation_in(reg_activation_7_11), .weight_in(reg_weight_6_12), .partial_sum_in(reg_psum_6_12), .reg_activation(reg_activation_7_12), .reg_weight(reg_weight_7_12), .reg_partial_sum(reg_psum_7_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_13( .activation_in(reg_activation_7_12), .weight_in(reg_weight_6_13), .partial_sum_in(reg_psum_6_13), .reg_activation(reg_activation_7_13), .reg_weight(reg_weight_7_13), .reg_partial_sum(reg_psum_7_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_14( .activation_in(reg_activation_7_13), .weight_in(reg_weight_6_14), .partial_sum_in(reg_psum_6_14), .reg_activation(reg_activation_7_14), .reg_weight(reg_weight_7_14), .reg_partial_sum(reg_psum_7_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_15( .activation_in(reg_activation_7_14), .weight_in(reg_weight_6_15), .partial_sum_in(reg_psum_6_15), .reg_activation(reg_activation_7_15), .reg_weight(reg_weight_7_15), .reg_partial_sum(reg_psum_7_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_16( .activation_in(reg_activation_7_15), .weight_in(reg_weight_6_16), .partial_sum_in(reg_psum_6_16), .reg_activation(reg_activation_7_16), .reg_weight(reg_weight_7_16), .reg_partial_sum(reg_psum_7_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_17( .activation_in(reg_activation_7_16), .weight_in(reg_weight_6_17), .partial_sum_in(reg_psum_6_17), .reg_activation(reg_activation_7_17), .reg_weight(reg_weight_7_17), .reg_partial_sum(reg_psum_7_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_18( .activation_in(reg_activation_7_17), .weight_in(reg_weight_6_18), .partial_sum_in(reg_psum_6_18), .reg_activation(reg_activation_7_18), .reg_weight(reg_weight_7_18), .reg_partial_sum(reg_psum_7_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_19( .activation_in(reg_activation_7_18), .weight_in(reg_weight_6_19), .partial_sum_in(reg_psum_6_19), .reg_activation(reg_activation_7_19), .reg_weight(reg_weight_7_19), .reg_partial_sum(reg_psum_7_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_20( .activation_in(reg_activation_7_19), .weight_in(reg_weight_6_20), .partial_sum_in(reg_psum_6_20), .reg_activation(reg_activation_7_20), .reg_weight(reg_weight_7_20), .reg_partial_sum(reg_psum_7_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_21( .activation_in(reg_activation_7_20), .weight_in(reg_weight_6_21), .partial_sum_in(reg_psum_6_21), .reg_activation(reg_activation_7_21), .reg_weight(reg_weight_7_21), .reg_partial_sum(reg_psum_7_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_22( .activation_in(reg_activation_7_21), .weight_in(reg_weight_6_22), .partial_sum_in(reg_psum_6_22), .reg_activation(reg_activation_7_22), .reg_weight(reg_weight_7_22), .reg_partial_sum(reg_psum_7_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_23( .activation_in(reg_activation_7_22), .weight_in(reg_weight_6_23), .partial_sum_in(reg_psum_6_23), .reg_activation(reg_activation_7_23), .reg_weight(reg_weight_7_23), .reg_partial_sum(reg_psum_7_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_24( .activation_in(reg_activation_7_23), .weight_in(reg_weight_6_24), .partial_sum_in(reg_psum_6_24), .reg_activation(reg_activation_7_24), .reg_weight(reg_weight_7_24), .reg_partial_sum(reg_psum_7_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_25( .activation_in(reg_activation_7_24), .weight_in(reg_weight_6_25), .partial_sum_in(reg_psum_6_25), .reg_activation(reg_activation_7_25), .reg_weight(reg_weight_7_25), .reg_partial_sum(reg_psum_7_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_26( .activation_in(reg_activation_7_25), .weight_in(reg_weight_6_26), .partial_sum_in(reg_psum_6_26), .reg_activation(reg_activation_7_26), .reg_weight(reg_weight_7_26), .reg_partial_sum(reg_psum_7_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_27( .activation_in(reg_activation_7_26), .weight_in(reg_weight_6_27), .partial_sum_in(reg_psum_6_27), .reg_activation(reg_activation_7_27), .reg_weight(reg_weight_7_27), .reg_partial_sum(reg_psum_7_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_28( .activation_in(reg_activation_7_27), .weight_in(reg_weight_6_28), .partial_sum_in(reg_psum_6_28), .reg_activation(reg_activation_7_28), .reg_weight(reg_weight_7_28), .reg_partial_sum(reg_psum_7_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_29( .activation_in(reg_activation_7_28), .weight_in(reg_weight_6_29), .partial_sum_in(reg_psum_6_29), .reg_activation(reg_activation_7_29), .reg_weight(reg_weight_7_29), .reg_partial_sum(reg_psum_7_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_30( .activation_in(reg_activation_7_29), .weight_in(reg_weight_6_30), .partial_sum_in(reg_psum_6_30), .reg_activation(reg_activation_7_30), .reg_weight(reg_weight_7_30), .reg_partial_sum(reg_psum_7_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_31( .activation_in(reg_activation_7_30), .weight_in(reg_weight_6_31), .partial_sum_in(reg_psum_6_31), .reg_activation(reg_activation_7_31), .reg_weight(reg_weight_7_31), .reg_partial_sum(reg_psum_7_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_32( .activation_in(reg_activation_7_31), .weight_in(reg_weight_6_32), .partial_sum_in(reg_psum_6_32), .reg_activation(reg_activation_7_32), .reg_weight(reg_weight_7_32), .reg_partial_sum(reg_psum_7_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_33( .activation_in(reg_activation_7_32), .weight_in(reg_weight_6_33), .partial_sum_in(reg_psum_6_33), .reg_activation(reg_activation_7_33), .reg_weight(reg_weight_7_33), .reg_partial_sum(reg_psum_7_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_34( .activation_in(reg_activation_7_33), .weight_in(reg_weight_6_34), .partial_sum_in(reg_psum_6_34), .reg_activation(reg_activation_7_34), .reg_weight(reg_weight_7_34), .reg_partial_sum(reg_psum_7_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_35( .activation_in(reg_activation_7_34), .weight_in(reg_weight_6_35), .partial_sum_in(reg_psum_6_35), .reg_activation(reg_activation_7_35), .reg_weight(reg_weight_7_35), .reg_partial_sum(reg_psum_7_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_36( .activation_in(reg_activation_7_35), .weight_in(reg_weight_6_36), .partial_sum_in(reg_psum_6_36), .reg_activation(reg_activation_7_36), .reg_weight(reg_weight_7_36), .reg_partial_sum(reg_psum_7_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_37( .activation_in(reg_activation_7_36), .weight_in(reg_weight_6_37), .partial_sum_in(reg_psum_6_37), .reg_activation(reg_activation_7_37), .reg_weight(reg_weight_7_37), .reg_partial_sum(reg_psum_7_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_38( .activation_in(reg_activation_7_37), .weight_in(reg_weight_6_38), .partial_sum_in(reg_psum_6_38), .reg_activation(reg_activation_7_38), .reg_weight(reg_weight_7_38), .reg_partial_sum(reg_psum_7_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_39( .activation_in(reg_activation_7_38), .weight_in(reg_weight_6_39), .partial_sum_in(reg_psum_6_39), .reg_activation(reg_activation_7_39), .reg_weight(reg_weight_7_39), .reg_partial_sum(reg_psum_7_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_40( .activation_in(reg_activation_7_39), .weight_in(reg_weight_6_40), .partial_sum_in(reg_psum_6_40), .reg_activation(reg_activation_7_40), .reg_weight(reg_weight_7_40), .reg_partial_sum(reg_psum_7_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_41( .activation_in(reg_activation_7_40), .weight_in(reg_weight_6_41), .partial_sum_in(reg_psum_6_41), .reg_activation(reg_activation_7_41), .reg_weight(reg_weight_7_41), .reg_partial_sum(reg_psum_7_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_42( .activation_in(reg_activation_7_41), .weight_in(reg_weight_6_42), .partial_sum_in(reg_psum_6_42), .reg_activation(reg_activation_7_42), .reg_weight(reg_weight_7_42), .reg_partial_sum(reg_psum_7_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_43( .activation_in(reg_activation_7_42), .weight_in(reg_weight_6_43), .partial_sum_in(reg_psum_6_43), .reg_activation(reg_activation_7_43), .reg_weight(reg_weight_7_43), .reg_partial_sum(reg_psum_7_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_44( .activation_in(reg_activation_7_43), .weight_in(reg_weight_6_44), .partial_sum_in(reg_psum_6_44), .reg_activation(reg_activation_7_44), .reg_weight(reg_weight_7_44), .reg_partial_sum(reg_psum_7_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_45( .activation_in(reg_activation_7_44), .weight_in(reg_weight_6_45), .partial_sum_in(reg_psum_6_45), .reg_activation(reg_activation_7_45), .reg_weight(reg_weight_7_45), .reg_partial_sum(reg_psum_7_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_46( .activation_in(reg_activation_7_45), .weight_in(reg_weight_6_46), .partial_sum_in(reg_psum_6_46), .reg_activation(reg_activation_7_46), .reg_weight(reg_weight_7_46), .reg_partial_sum(reg_psum_7_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_47( .activation_in(reg_activation_7_46), .weight_in(reg_weight_6_47), .partial_sum_in(reg_psum_6_47), .reg_activation(reg_activation_7_47), .reg_weight(reg_weight_7_47), .reg_partial_sum(reg_psum_7_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_48( .activation_in(reg_activation_7_47), .weight_in(reg_weight_6_48), .partial_sum_in(reg_psum_6_48), .reg_activation(reg_activation_7_48), .reg_weight(reg_weight_7_48), .reg_partial_sum(reg_psum_7_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_49( .activation_in(reg_activation_7_48), .weight_in(reg_weight_6_49), .partial_sum_in(reg_psum_6_49), .reg_activation(reg_activation_7_49), .reg_weight(reg_weight_7_49), .reg_partial_sum(reg_psum_7_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_50( .activation_in(reg_activation_7_49), .weight_in(reg_weight_6_50), .partial_sum_in(reg_psum_6_50), .reg_activation(reg_activation_7_50), .reg_weight(reg_weight_7_50), .reg_partial_sum(reg_psum_7_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_51( .activation_in(reg_activation_7_50), .weight_in(reg_weight_6_51), .partial_sum_in(reg_psum_6_51), .reg_activation(reg_activation_7_51), .reg_weight(reg_weight_7_51), .reg_partial_sum(reg_psum_7_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_52( .activation_in(reg_activation_7_51), .weight_in(reg_weight_6_52), .partial_sum_in(reg_psum_6_52), .reg_activation(reg_activation_7_52), .reg_weight(reg_weight_7_52), .reg_partial_sum(reg_psum_7_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_53( .activation_in(reg_activation_7_52), .weight_in(reg_weight_6_53), .partial_sum_in(reg_psum_6_53), .reg_activation(reg_activation_7_53), .reg_weight(reg_weight_7_53), .reg_partial_sum(reg_psum_7_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_54( .activation_in(reg_activation_7_53), .weight_in(reg_weight_6_54), .partial_sum_in(reg_psum_6_54), .reg_activation(reg_activation_7_54), .reg_weight(reg_weight_7_54), .reg_partial_sum(reg_psum_7_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_55( .activation_in(reg_activation_7_54), .weight_in(reg_weight_6_55), .partial_sum_in(reg_psum_6_55), .reg_activation(reg_activation_7_55), .reg_weight(reg_weight_7_55), .reg_partial_sum(reg_psum_7_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_56( .activation_in(reg_activation_7_55), .weight_in(reg_weight_6_56), .partial_sum_in(reg_psum_6_56), .reg_activation(reg_activation_7_56), .reg_weight(reg_weight_7_56), .reg_partial_sum(reg_psum_7_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_57( .activation_in(reg_activation_7_56), .weight_in(reg_weight_6_57), .partial_sum_in(reg_psum_6_57), .reg_activation(reg_activation_7_57), .reg_weight(reg_weight_7_57), .reg_partial_sum(reg_psum_7_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_58( .activation_in(reg_activation_7_57), .weight_in(reg_weight_6_58), .partial_sum_in(reg_psum_6_58), .reg_activation(reg_activation_7_58), .reg_weight(reg_weight_7_58), .reg_partial_sum(reg_psum_7_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_59( .activation_in(reg_activation_7_58), .weight_in(reg_weight_6_59), .partial_sum_in(reg_psum_6_59), .reg_activation(reg_activation_7_59), .reg_weight(reg_weight_7_59), .reg_partial_sum(reg_psum_7_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_60( .activation_in(reg_activation_7_59), .weight_in(reg_weight_6_60), .partial_sum_in(reg_psum_6_60), .reg_activation(reg_activation_7_60), .reg_weight(reg_weight_7_60), .reg_partial_sum(reg_psum_7_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_61( .activation_in(reg_activation_7_60), .weight_in(reg_weight_6_61), .partial_sum_in(reg_psum_6_61), .reg_activation(reg_activation_7_61), .reg_weight(reg_weight_7_61), .reg_partial_sum(reg_psum_7_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_62( .activation_in(reg_activation_7_61), .weight_in(reg_weight_6_62), .partial_sum_in(reg_psum_6_62), .reg_activation(reg_activation_7_62), .reg_weight(reg_weight_7_62), .reg_partial_sum(reg_psum_7_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_63( .activation_in(reg_activation_7_62), .weight_in(reg_weight_6_63), .partial_sum_in(reg_psum_6_63), .reg_weight(reg_weight_7_63), .reg_partial_sum(reg_psum_7_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_0( .activation_in(in_activation_8), .weight_in(reg_weight_7_0), .partial_sum_in(reg_psum_7_0), .reg_activation(reg_activation_8_0), .reg_weight(reg_weight_8_0), .reg_partial_sum(reg_psum_8_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_1( .activation_in(reg_activation_8_0), .weight_in(reg_weight_7_1), .partial_sum_in(reg_psum_7_1), .reg_activation(reg_activation_8_1), .reg_weight(reg_weight_8_1), .reg_partial_sum(reg_psum_8_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_2( .activation_in(reg_activation_8_1), .weight_in(reg_weight_7_2), .partial_sum_in(reg_psum_7_2), .reg_activation(reg_activation_8_2), .reg_weight(reg_weight_8_2), .reg_partial_sum(reg_psum_8_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_3( .activation_in(reg_activation_8_2), .weight_in(reg_weight_7_3), .partial_sum_in(reg_psum_7_3), .reg_activation(reg_activation_8_3), .reg_weight(reg_weight_8_3), .reg_partial_sum(reg_psum_8_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_4( .activation_in(reg_activation_8_3), .weight_in(reg_weight_7_4), .partial_sum_in(reg_psum_7_4), .reg_activation(reg_activation_8_4), .reg_weight(reg_weight_8_4), .reg_partial_sum(reg_psum_8_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_5( .activation_in(reg_activation_8_4), .weight_in(reg_weight_7_5), .partial_sum_in(reg_psum_7_5), .reg_activation(reg_activation_8_5), .reg_weight(reg_weight_8_5), .reg_partial_sum(reg_psum_8_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_6( .activation_in(reg_activation_8_5), .weight_in(reg_weight_7_6), .partial_sum_in(reg_psum_7_6), .reg_activation(reg_activation_8_6), .reg_weight(reg_weight_8_6), .reg_partial_sum(reg_psum_8_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_7( .activation_in(reg_activation_8_6), .weight_in(reg_weight_7_7), .partial_sum_in(reg_psum_7_7), .reg_activation(reg_activation_8_7), .reg_weight(reg_weight_8_7), .reg_partial_sum(reg_psum_8_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_8( .activation_in(reg_activation_8_7), .weight_in(reg_weight_7_8), .partial_sum_in(reg_psum_7_8), .reg_activation(reg_activation_8_8), .reg_weight(reg_weight_8_8), .reg_partial_sum(reg_psum_8_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_9( .activation_in(reg_activation_8_8), .weight_in(reg_weight_7_9), .partial_sum_in(reg_psum_7_9), .reg_activation(reg_activation_8_9), .reg_weight(reg_weight_8_9), .reg_partial_sum(reg_psum_8_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_10( .activation_in(reg_activation_8_9), .weight_in(reg_weight_7_10), .partial_sum_in(reg_psum_7_10), .reg_activation(reg_activation_8_10), .reg_weight(reg_weight_8_10), .reg_partial_sum(reg_psum_8_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_11( .activation_in(reg_activation_8_10), .weight_in(reg_weight_7_11), .partial_sum_in(reg_psum_7_11), .reg_activation(reg_activation_8_11), .reg_weight(reg_weight_8_11), .reg_partial_sum(reg_psum_8_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_12( .activation_in(reg_activation_8_11), .weight_in(reg_weight_7_12), .partial_sum_in(reg_psum_7_12), .reg_activation(reg_activation_8_12), .reg_weight(reg_weight_8_12), .reg_partial_sum(reg_psum_8_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_13( .activation_in(reg_activation_8_12), .weight_in(reg_weight_7_13), .partial_sum_in(reg_psum_7_13), .reg_activation(reg_activation_8_13), .reg_weight(reg_weight_8_13), .reg_partial_sum(reg_psum_8_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_14( .activation_in(reg_activation_8_13), .weight_in(reg_weight_7_14), .partial_sum_in(reg_psum_7_14), .reg_activation(reg_activation_8_14), .reg_weight(reg_weight_8_14), .reg_partial_sum(reg_psum_8_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_15( .activation_in(reg_activation_8_14), .weight_in(reg_weight_7_15), .partial_sum_in(reg_psum_7_15), .reg_activation(reg_activation_8_15), .reg_weight(reg_weight_8_15), .reg_partial_sum(reg_psum_8_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_16( .activation_in(reg_activation_8_15), .weight_in(reg_weight_7_16), .partial_sum_in(reg_psum_7_16), .reg_activation(reg_activation_8_16), .reg_weight(reg_weight_8_16), .reg_partial_sum(reg_psum_8_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_17( .activation_in(reg_activation_8_16), .weight_in(reg_weight_7_17), .partial_sum_in(reg_psum_7_17), .reg_activation(reg_activation_8_17), .reg_weight(reg_weight_8_17), .reg_partial_sum(reg_psum_8_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_18( .activation_in(reg_activation_8_17), .weight_in(reg_weight_7_18), .partial_sum_in(reg_psum_7_18), .reg_activation(reg_activation_8_18), .reg_weight(reg_weight_8_18), .reg_partial_sum(reg_psum_8_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_19( .activation_in(reg_activation_8_18), .weight_in(reg_weight_7_19), .partial_sum_in(reg_psum_7_19), .reg_activation(reg_activation_8_19), .reg_weight(reg_weight_8_19), .reg_partial_sum(reg_psum_8_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_20( .activation_in(reg_activation_8_19), .weight_in(reg_weight_7_20), .partial_sum_in(reg_psum_7_20), .reg_activation(reg_activation_8_20), .reg_weight(reg_weight_8_20), .reg_partial_sum(reg_psum_8_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_21( .activation_in(reg_activation_8_20), .weight_in(reg_weight_7_21), .partial_sum_in(reg_psum_7_21), .reg_activation(reg_activation_8_21), .reg_weight(reg_weight_8_21), .reg_partial_sum(reg_psum_8_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_22( .activation_in(reg_activation_8_21), .weight_in(reg_weight_7_22), .partial_sum_in(reg_psum_7_22), .reg_activation(reg_activation_8_22), .reg_weight(reg_weight_8_22), .reg_partial_sum(reg_psum_8_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_23( .activation_in(reg_activation_8_22), .weight_in(reg_weight_7_23), .partial_sum_in(reg_psum_7_23), .reg_activation(reg_activation_8_23), .reg_weight(reg_weight_8_23), .reg_partial_sum(reg_psum_8_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_24( .activation_in(reg_activation_8_23), .weight_in(reg_weight_7_24), .partial_sum_in(reg_psum_7_24), .reg_activation(reg_activation_8_24), .reg_weight(reg_weight_8_24), .reg_partial_sum(reg_psum_8_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_25( .activation_in(reg_activation_8_24), .weight_in(reg_weight_7_25), .partial_sum_in(reg_psum_7_25), .reg_activation(reg_activation_8_25), .reg_weight(reg_weight_8_25), .reg_partial_sum(reg_psum_8_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_26( .activation_in(reg_activation_8_25), .weight_in(reg_weight_7_26), .partial_sum_in(reg_psum_7_26), .reg_activation(reg_activation_8_26), .reg_weight(reg_weight_8_26), .reg_partial_sum(reg_psum_8_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_27( .activation_in(reg_activation_8_26), .weight_in(reg_weight_7_27), .partial_sum_in(reg_psum_7_27), .reg_activation(reg_activation_8_27), .reg_weight(reg_weight_8_27), .reg_partial_sum(reg_psum_8_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_28( .activation_in(reg_activation_8_27), .weight_in(reg_weight_7_28), .partial_sum_in(reg_psum_7_28), .reg_activation(reg_activation_8_28), .reg_weight(reg_weight_8_28), .reg_partial_sum(reg_psum_8_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_29( .activation_in(reg_activation_8_28), .weight_in(reg_weight_7_29), .partial_sum_in(reg_psum_7_29), .reg_activation(reg_activation_8_29), .reg_weight(reg_weight_8_29), .reg_partial_sum(reg_psum_8_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_30( .activation_in(reg_activation_8_29), .weight_in(reg_weight_7_30), .partial_sum_in(reg_psum_7_30), .reg_activation(reg_activation_8_30), .reg_weight(reg_weight_8_30), .reg_partial_sum(reg_psum_8_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_31( .activation_in(reg_activation_8_30), .weight_in(reg_weight_7_31), .partial_sum_in(reg_psum_7_31), .reg_activation(reg_activation_8_31), .reg_weight(reg_weight_8_31), .reg_partial_sum(reg_psum_8_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_32( .activation_in(reg_activation_8_31), .weight_in(reg_weight_7_32), .partial_sum_in(reg_psum_7_32), .reg_activation(reg_activation_8_32), .reg_weight(reg_weight_8_32), .reg_partial_sum(reg_psum_8_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_33( .activation_in(reg_activation_8_32), .weight_in(reg_weight_7_33), .partial_sum_in(reg_psum_7_33), .reg_activation(reg_activation_8_33), .reg_weight(reg_weight_8_33), .reg_partial_sum(reg_psum_8_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_34( .activation_in(reg_activation_8_33), .weight_in(reg_weight_7_34), .partial_sum_in(reg_psum_7_34), .reg_activation(reg_activation_8_34), .reg_weight(reg_weight_8_34), .reg_partial_sum(reg_psum_8_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_35( .activation_in(reg_activation_8_34), .weight_in(reg_weight_7_35), .partial_sum_in(reg_psum_7_35), .reg_activation(reg_activation_8_35), .reg_weight(reg_weight_8_35), .reg_partial_sum(reg_psum_8_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_36( .activation_in(reg_activation_8_35), .weight_in(reg_weight_7_36), .partial_sum_in(reg_psum_7_36), .reg_activation(reg_activation_8_36), .reg_weight(reg_weight_8_36), .reg_partial_sum(reg_psum_8_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_37( .activation_in(reg_activation_8_36), .weight_in(reg_weight_7_37), .partial_sum_in(reg_psum_7_37), .reg_activation(reg_activation_8_37), .reg_weight(reg_weight_8_37), .reg_partial_sum(reg_psum_8_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_38( .activation_in(reg_activation_8_37), .weight_in(reg_weight_7_38), .partial_sum_in(reg_psum_7_38), .reg_activation(reg_activation_8_38), .reg_weight(reg_weight_8_38), .reg_partial_sum(reg_psum_8_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_39( .activation_in(reg_activation_8_38), .weight_in(reg_weight_7_39), .partial_sum_in(reg_psum_7_39), .reg_activation(reg_activation_8_39), .reg_weight(reg_weight_8_39), .reg_partial_sum(reg_psum_8_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_40( .activation_in(reg_activation_8_39), .weight_in(reg_weight_7_40), .partial_sum_in(reg_psum_7_40), .reg_activation(reg_activation_8_40), .reg_weight(reg_weight_8_40), .reg_partial_sum(reg_psum_8_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_41( .activation_in(reg_activation_8_40), .weight_in(reg_weight_7_41), .partial_sum_in(reg_psum_7_41), .reg_activation(reg_activation_8_41), .reg_weight(reg_weight_8_41), .reg_partial_sum(reg_psum_8_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_42( .activation_in(reg_activation_8_41), .weight_in(reg_weight_7_42), .partial_sum_in(reg_psum_7_42), .reg_activation(reg_activation_8_42), .reg_weight(reg_weight_8_42), .reg_partial_sum(reg_psum_8_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_43( .activation_in(reg_activation_8_42), .weight_in(reg_weight_7_43), .partial_sum_in(reg_psum_7_43), .reg_activation(reg_activation_8_43), .reg_weight(reg_weight_8_43), .reg_partial_sum(reg_psum_8_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_44( .activation_in(reg_activation_8_43), .weight_in(reg_weight_7_44), .partial_sum_in(reg_psum_7_44), .reg_activation(reg_activation_8_44), .reg_weight(reg_weight_8_44), .reg_partial_sum(reg_psum_8_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_45( .activation_in(reg_activation_8_44), .weight_in(reg_weight_7_45), .partial_sum_in(reg_psum_7_45), .reg_activation(reg_activation_8_45), .reg_weight(reg_weight_8_45), .reg_partial_sum(reg_psum_8_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_46( .activation_in(reg_activation_8_45), .weight_in(reg_weight_7_46), .partial_sum_in(reg_psum_7_46), .reg_activation(reg_activation_8_46), .reg_weight(reg_weight_8_46), .reg_partial_sum(reg_psum_8_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_47( .activation_in(reg_activation_8_46), .weight_in(reg_weight_7_47), .partial_sum_in(reg_psum_7_47), .reg_activation(reg_activation_8_47), .reg_weight(reg_weight_8_47), .reg_partial_sum(reg_psum_8_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_48( .activation_in(reg_activation_8_47), .weight_in(reg_weight_7_48), .partial_sum_in(reg_psum_7_48), .reg_activation(reg_activation_8_48), .reg_weight(reg_weight_8_48), .reg_partial_sum(reg_psum_8_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_49( .activation_in(reg_activation_8_48), .weight_in(reg_weight_7_49), .partial_sum_in(reg_psum_7_49), .reg_activation(reg_activation_8_49), .reg_weight(reg_weight_8_49), .reg_partial_sum(reg_psum_8_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_50( .activation_in(reg_activation_8_49), .weight_in(reg_weight_7_50), .partial_sum_in(reg_psum_7_50), .reg_activation(reg_activation_8_50), .reg_weight(reg_weight_8_50), .reg_partial_sum(reg_psum_8_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_51( .activation_in(reg_activation_8_50), .weight_in(reg_weight_7_51), .partial_sum_in(reg_psum_7_51), .reg_activation(reg_activation_8_51), .reg_weight(reg_weight_8_51), .reg_partial_sum(reg_psum_8_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_52( .activation_in(reg_activation_8_51), .weight_in(reg_weight_7_52), .partial_sum_in(reg_psum_7_52), .reg_activation(reg_activation_8_52), .reg_weight(reg_weight_8_52), .reg_partial_sum(reg_psum_8_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_53( .activation_in(reg_activation_8_52), .weight_in(reg_weight_7_53), .partial_sum_in(reg_psum_7_53), .reg_activation(reg_activation_8_53), .reg_weight(reg_weight_8_53), .reg_partial_sum(reg_psum_8_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_54( .activation_in(reg_activation_8_53), .weight_in(reg_weight_7_54), .partial_sum_in(reg_psum_7_54), .reg_activation(reg_activation_8_54), .reg_weight(reg_weight_8_54), .reg_partial_sum(reg_psum_8_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_55( .activation_in(reg_activation_8_54), .weight_in(reg_weight_7_55), .partial_sum_in(reg_psum_7_55), .reg_activation(reg_activation_8_55), .reg_weight(reg_weight_8_55), .reg_partial_sum(reg_psum_8_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_56( .activation_in(reg_activation_8_55), .weight_in(reg_weight_7_56), .partial_sum_in(reg_psum_7_56), .reg_activation(reg_activation_8_56), .reg_weight(reg_weight_8_56), .reg_partial_sum(reg_psum_8_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_57( .activation_in(reg_activation_8_56), .weight_in(reg_weight_7_57), .partial_sum_in(reg_psum_7_57), .reg_activation(reg_activation_8_57), .reg_weight(reg_weight_8_57), .reg_partial_sum(reg_psum_8_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_58( .activation_in(reg_activation_8_57), .weight_in(reg_weight_7_58), .partial_sum_in(reg_psum_7_58), .reg_activation(reg_activation_8_58), .reg_weight(reg_weight_8_58), .reg_partial_sum(reg_psum_8_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_59( .activation_in(reg_activation_8_58), .weight_in(reg_weight_7_59), .partial_sum_in(reg_psum_7_59), .reg_activation(reg_activation_8_59), .reg_weight(reg_weight_8_59), .reg_partial_sum(reg_psum_8_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_60( .activation_in(reg_activation_8_59), .weight_in(reg_weight_7_60), .partial_sum_in(reg_psum_7_60), .reg_activation(reg_activation_8_60), .reg_weight(reg_weight_8_60), .reg_partial_sum(reg_psum_8_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_61( .activation_in(reg_activation_8_60), .weight_in(reg_weight_7_61), .partial_sum_in(reg_psum_7_61), .reg_activation(reg_activation_8_61), .reg_weight(reg_weight_8_61), .reg_partial_sum(reg_psum_8_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_62( .activation_in(reg_activation_8_61), .weight_in(reg_weight_7_62), .partial_sum_in(reg_psum_7_62), .reg_activation(reg_activation_8_62), .reg_weight(reg_weight_8_62), .reg_partial_sum(reg_psum_8_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_63( .activation_in(reg_activation_8_62), .weight_in(reg_weight_7_63), .partial_sum_in(reg_psum_7_63), .reg_weight(reg_weight_8_63), .reg_partial_sum(reg_psum_8_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_0( .activation_in(in_activation_9), .weight_in(reg_weight_8_0), .partial_sum_in(reg_psum_8_0), .reg_activation(reg_activation_9_0), .reg_weight(reg_weight_9_0), .reg_partial_sum(reg_psum_9_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_1( .activation_in(reg_activation_9_0), .weight_in(reg_weight_8_1), .partial_sum_in(reg_psum_8_1), .reg_activation(reg_activation_9_1), .reg_weight(reg_weight_9_1), .reg_partial_sum(reg_psum_9_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_2( .activation_in(reg_activation_9_1), .weight_in(reg_weight_8_2), .partial_sum_in(reg_psum_8_2), .reg_activation(reg_activation_9_2), .reg_weight(reg_weight_9_2), .reg_partial_sum(reg_psum_9_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_3( .activation_in(reg_activation_9_2), .weight_in(reg_weight_8_3), .partial_sum_in(reg_psum_8_3), .reg_activation(reg_activation_9_3), .reg_weight(reg_weight_9_3), .reg_partial_sum(reg_psum_9_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_4( .activation_in(reg_activation_9_3), .weight_in(reg_weight_8_4), .partial_sum_in(reg_psum_8_4), .reg_activation(reg_activation_9_4), .reg_weight(reg_weight_9_4), .reg_partial_sum(reg_psum_9_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_5( .activation_in(reg_activation_9_4), .weight_in(reg_weight_8_5), .partial_sum_in(reg_psum_8_5), .reg_activation(reg_activation_9_5), .reg_weight(reg_weight_9_5), .reg_partial_sum(reg_psum_9_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_6( .activation_in(reg_activation_9_5), .weight_in(reg_weight_8_6), .partial_sum_in(reg_psum_8_6), .reg_activation(reg_activation_9_6), .reg_weight(reg_weight_9_6), .reg_partial_sum(reg_psum_9_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_7( .activation_in(reg_activation_9_6), .weight_in(reg_weight_8_7), .partial_sum_in(reg_psum_8_7), .reg_activation(reg_activation_9_7), .reg_weight(reg_weight_9_7), .reg_partial_sum(reg_psum_9_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_8( .activation_in(reg_activation_9_7), .weight_in(reg_weight_8_8), .partial_sum_in(reg_psum_8_8), .reg_activation(reg_activation_9_8), .reg_weight(reg_weight_9_8), .reg_partial_sum(reg_psum_9_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_9( .activation_in(reg_activation_9_8), .weight_in(reg_weight_8_9), .partial_sum_in(reg_psum_8_9), .reg_activation(reg_activation_9_9), .reg_weight(reg_weight_9_9), .reg_partial_sum(reg_psum_9_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_10( .activation_in(reg_activation_9_9), .weight_in(reg_weight_8_10), .partial_sum_in(reg_psum_8_10), .reg_activation(reg_activation_9_10), .reg_weight(reg_weight_9_10), .reg_partial_sum(reg_psum_9_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_11( .activation_in(reg_activation_9_10), .weight_in(reg_weight_8_11), .partial_sum_in(reg_psum_8_11), .reg_activation(reg_activation_9_11), .reg_weight(reg_weight_9_11), .reg_partial_sum(reg_psum_9_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_12( .activation_in(reg_activation_9_11), .weight_in(reg_weight_8_12), .partial_sum_in(reg_psum_8_12), .reg_activation(reg_activation_9_12), .reg_weight(reg_weight_9_12), .reg_partial_sum(reg_psum_9_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_13( .activation_in(reg_activation_9_12), .weight_in(reg_weight_8_13), .partial_sum_in(reg_psum_8_13), .reg_activation(reg_activation_9_13), .reg_weight(reg_weight_9_13), .reg_partial_sum(reg_psum_9_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_14( .activation_in(reg_activation_9_13), .weight_in(reg_weight_8_14), .partial_sum_in(reg_psum_8_14), .reg_activation(reg_activation_9_14), .reg_weight(reg_weight_9_14), .reg_partial_sum(reg_psum_9_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_15( .activation_in(reg_activation_9_14), .weight_in(reg_weight_8_15), .partial_sum_in(reg_psum_8_15), .reg_activation(reg_activation_9_15), .reg_weight(reg_weight_9_15), .reg_partial_sum(reg_psum_9_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_16( .activation_in(reg_activation_9_15), .weight_in(reg_weight_8_16), .partial_sum_in(reg_psum_8_16), .reg_activation(reg_activation_9_16), .reg_weight(reg_weight_9_16), .reg_partial_sum(reg_psum_9_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_17( .activation_in(reg_activation_9_16), .weight_in(reg_weight_8_17), .partial_sum_in(reg_psum_8_17), .reg_activation(reg_activation_9_17), .reg_weight(reg_weight_9_17), .reg_partial_sum(reg_psum_9_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_18( .activation_in(reg_activation_9_17), .weight_in(reg_weight_8_18), .partial_sum_in(reg_psum_8_18), .reg_activation(reg_activation_9_18), .reg_weight(reg_weight_9_18), .reg_partial_sum(reg_psum_9_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_19( .activation_in(reg_activation_9_18), .weight_in(reg_weight_8_19), .partial_sum_in(reg_psum_8_19), .reg_activation(reg_activation_9_19), .reg_weight(reg_weight_9_19), .reg_partial_sum(reg_psum_9_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_20( .activation_in(reg_activation_9_19), .weight_in(reg_weight_8_20), .partial_sum_in(reg_psum_8_20), .reg_activation(reg_activation_9_20), .reg_weight(reg_weight_9_20), .reg_partial_sum(reg_psum_9_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_21( .activation_in(reg_activation_9_20), .weight_in(reg_weight_8_21), .partial_sum_in(reg_psum_8_21), .reg_activation(reg_activation_9_21), .reg_weight(reg_weight_9_21), .reg_partial_sum(reg_psum_9_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_22( .activation_in(reg_activation_9_21), .weight_in(reg_weight_8_22), .partial_sum_in(reg_psum_8_22), .reg_activation(reg_activation_9_22), .reg_weight(reg_weight_9_22), .reg_partial_sum(reg_psum_9_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_23( .activation_in(reg_activation_9_22), .weight_in(reg_weight_8_23), .partial_sum_in(reg_psum_8_23), .reg_activation(reg_activation_9_23), .reg_weight(reg_weight_9_23), .reg_partial_sum(reg_psum_9_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_24( .activation_in(reg_activation_9_23), .weight_in(reg_weight_8_24), .partial_sum_in(reg_psum_8_24), .reg_activation(reg_activation_9_24), .reg_weight(reg_weight_9_24), .reg_partial_sum(reg_psum_9_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_25( .activation_in(reg_activation_9_24), .weight_in(reg_weight_8_25), .partial_sum_in(reg_psum_8_25), .reg_activation(reg_activation_9_25), .reg_weight(reg_weight_9_25), .reg_partial_sum(reg_psum_9_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_26( .activation_in(reg_activation_9_25), .weight_in(reg_weight_8_26), .partial_sum_in(reg_psum_8_26), .reg_activation(reg_activation_9_26), .reg_weight(reg_weight_9_26), .reg_partial_sum(reg_psum_9_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_27( .activation_in(reg_activation_9_26), .weight_in(reg_weight_8_27), .partial_sum_in(reg_psum_8_27), .reg_activation(reg_activation_9_27), .reg_weight(reg_weight_9_27), .reg_partial_sum(reg_psum_9_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_28( .activation_in(reg_activation_9_27), .weight_in(reg_weight_8_28), .partial_sum_in(reg_psum_8_28), .reg_activation(reg_activation_9_28), .reg_weight(reg_weight_9_28), .reg_partial_sum(reg_psum_9_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_29( .activation_in(reg_activation_9_28), .weight_in(reg_weight_8_29), .partial_sum_in(reg_psum_8_29), .reg_activation(reg_activation_9_29), .reg_weight(reg_weight_9_29), .reg_partial_sum(reg_psum_9_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_30( .activation_in(reg_activation_9_29), .weight_in(reg_weight_8_30), .partial_sum_in(reg_psum_8_30), .reg_activation(reg_activation_9_30), .reg_weight(reg_weight_9_30), .reg_partial_sum(reg_psum_9_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_31( .activation_in(reg_activation_9_30), .weight_in(reg_weight_8_31), .partial_sum_in(reg_psum_8_31), .reg_activation(reg_activation_9_31), .reg_weight(reg_weight_9_31), .reg_partial_sum(reg_psum_9_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_32( .activation_in(reg_activation_9_31), .weight_in(reg_weight_8_32), .partial_sum_in(reg_psum_8_32), .reg_activation(reg_activation_9_32), .reg_weight(reg_weight_9_32), .reg_partial_sum(reg_psum_9_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_33( .activation_in(reg_activation_9_32), .weight_in(reg_weight_8_33), .partial_sum_in(reg_psum_8_33), .reg_activation(reg_activation_9_33), .reg_weight(reg_weight_9_33), .reg_partial_sum(reg_psum_9_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_34( .activation_in(reg_activation_9_33), .weight_in(reg_weight_8_34), .partial_sum_in(reg_psum_8_34), .reg_activation(reg_activation_9_34), .reg_weight(reg_weight_9_34), .reg_partial_sum(reg_psum_9_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_35( .activation_in(reg_activation_9_34), .weight_in(reg_weight_8_35), .partial_sum_in(reg_psum_8_35), .reg_activation(reg_activation_9_35), .reg_weight(reg_weight_9_35), .reg_partial_sum(reg_psum_9_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_36( .activation_in(reg_activation_9_35), .weight_in(reg_weight_8_36), .partial_sum_in(reg_psum_8_36), .reg_activation(reg_activation_9_36), .reg_weight(reg_weight_9_36), .reg_partial_sum(reg_psum_9_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_37( .activation_in(reg_activation_9_36), .weight_in(reg_weight_8_37), .partial_sum_in(reg_psum_8_37), .reg_activation(reg_activation_9_37), .reg_weight(reg_weight_9_37), .reg_partial_sum(reg_psum_9_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_38( .activation_in(reg_activation_9_37), .weight_in(reg_weight_8_38), .partial_sum_in(reg_psum_8_38), .reg_activation(reg_activation_9_38), .reg_weight(reg_weight_9_38), .reg_partial_sum(reg_psum_9_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_39( .activation_in(reg_activation_9_38), .weight_in(reg_weight_8_39), .partial_sum_in(reg_psum_8_39), .reg_activation(reg_activation_9_39), .reg_weight(reg_weight_9_39), .reg_partial_sum(reg_psum_9_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_40( .activation_in(reg_activation_9_39), .weight_in(reg_weight_8_40), .partial_sum_in(reg_psum_8_40), .reg_activation(reg_activation_9_40), .reg_weight(reg_weight_9_40), .reg_partial_sum(reg_psum_9_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_41( .activation_in(reg_activation_9_40), .weight_in(reg_weight_8_41), .partial_sum_in(reg_psum_8_41), .reg_activation(reg_activation_9_41), .reg_weight(reg_weight_9_41), .reg_partial_sum(reg_psum_9_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_42( .activation_in(reg_activation_9_41), .weight_in(reg_weight_8_42), .partial_sum_in(reg_psum_8_42), .reg_activation(reg_activation_9_42), .reg_weight(reg_weight_9_42), .reg_partial_sum(reg_psum_9_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_43( .activation_in(reg_activation_9_42), .weight_in(reg_weight_8_43), .partial_sum_in(reg_psum_8_43), .reg_activation(reg_activation_9_43), .reg_weight(reg_weight_9_43), .reg_partial_sum(reg_psum_9_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_44( .activation_in(reg_activation_9_43), .weight_in(reg_weight_8_44), .partial_sum_in(reg_psum_8_44), .reg_activation(reg_activation_9_44), .reg_weight(reg_weight_9_44), .reg_partial_sum(reg_psum_9_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_45( .activation_in(reg_activation_9_44), .weight_in(reg_weight_8_45), .partial_sum_in(reg_psum_8_45), .reg_activation(reg_activation_9_45), .reg_weight(reg_weight_9_45), .reg_partial_sum(reg_psum_9_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_46( .activation_in(reg_activation_9_45), .weight_in(reg_weight_8_46), .partial_sum_in(reg_psum_8_46), .reg_activation(reg_activation_9_46), .reg_weight(reg_weight_9_46), .reg_partial_sum(reg_psum_9_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_47( .activation_in(reg_activation_9_46), .weight_in(reg_weight_8_47), .partial_sum_in(reg_psum_8_47), .reg_activation(reg_activation_9_47), .reg_weight(reg_weight_9_47), .reg_partial_sum(reg_psum_9_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_48( .activation_in(reg_activation_9_47), .weight_in(reg_weight_8_48), .partial_sum_in(reg_psum_8_48), .reg_activation(reg_activation_9_48), .reg_weight(reg_weight_9_48), .reg_partial_sum(reg_psum_9_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_49( .activation_in(reg_activation_9_48), .weight_in(reg_weight_8_49), .partial_sum_in(reg_psum_8_49), .reg_activation(reg_activation_9_49), .reg_weight(reg_weight_9_49), .reg_partial_sum(reg_psum_9_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_50( .activation_in(reg_activation_9_49), .weight_in(reg_weight_8_50), .partial_sum_in(reg_psum_8_50), .reg_activation(reg_activation_9_50), .reg_weight(reg_weight_9_50), .reg_partial_sum(reg_psum_9_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_51( .activation_in(reg_activation_9_50), .weight_in(reg_weight_8_51), .partial_sum_in(reg_psum_8_51), .reg_activation(reg_activation_9_51), .reg_weight(reg_weight_9_51), .reg_partial_sum(reg_psum_9_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_52( .activation_in(reg_activation_9_51), .weight_in(reg_weight_8_52), .partial_sum_in(reg_psum_8_52), .reg_activation(reg_activation_9_52), .reg_weight(reg_weight_9_52), .reg_partial_sum(reg_psum_9_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_53( .activation_in(reg_activation_9_52), .weight_in(reg_weight_8_53), .partial_sum_in(reg_psum_8_53), .reg_activation(reg_activation_9_53), .reg_weight(reg_weight_9_53), .reg_partial_sum(reg_psum_9_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_54( .activation_in(reg_activation_9_53), .weight_in(reg_weight_8_54), .partial_sum_in(reg_psum_8_54), .reg_activation(reg_activation_9_54), .reg_weight(reg_weight_9_54), .reg_partial_sum(reg_psum_9_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_55( .activation_in(reg_activation_9_54), .weight_in(reg_weight_8_55), .partial_sum_in(reg_psum_8_55), .reg_activation(reg_activation_9_55), .reg_weight(reg_weight_9_55), .reg_partial_sum(reg_psum_9_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_56( .activation_in(reg_activation_9_55), .weight_in(reg_weight_8_56), .partial_sum_in(reg_psum_8_56), .reg_activation(reg_activation_9_56), .reg_weight(reg_weight_9_56), .reg_partial_sum(reg_psum_9_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_57( .activation_in(reg_activation_9_56), .weight_in(reg_weight_8_57), .partial_sum_in(reg_psum_8_57), .reg_activation(reg_activation_9_57), .reg_weight(reg_weight_9_57), .reg_partial_sum(reg_psum_9_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_58( .activation_in(reg_activation_9_57), .weight_in(reg_weight_8_58), .partial_sum_in(reg_psum_8_58), .reg_activation(reg_activation_9_58), .reg_weight(reg_weight_9_58), .reg_partial_sum(reg_psum_9_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_59( .activation_in(reg_activation_9_58), .weight_in(reg_weight_8_59), .partial_sum_in(reg_psum_8_59), .reg_activation(reg_activation_9_59), .reg_weight(reg_weight_9_59), .reg_partial_sum(reg_psum_9_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_60( .activation_in(reg_activation_9_59), .weight_in(reg_weight_8_60), .partial_sum_in(reg_psum_8_60), .reg_activation(reg_activation_9_60), .reg_weight(reg_weight_9_60), .reg_partial_sum(reg_psum_9_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_61( .activation_in(reg_activation_9_60), .weight_in(reg_weight_8_61), .partial_sum_in(reg_psum_8_61), .reg_activation(reg_activation_9_61), .reg_weight(reg_weight_9_61), .reg_partial_sum(reg_psum_9_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_62( .activation_in(reg_activation_9_61), .weight_in(reg_weight_8_62), .partial_sum_in(reg_psum_8_62), .reg_activation(reg_activation_9_62), .reg_weight(reg_weight_9_62), .reg_partial_sum(reg_psum_9_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_63( .activation_in(reg_activation_9_62), .weight_in(reg_weight_8_63), .partial_sum_in(reg_psum_8_63), .reg_weight(reg_weight_9_63), .reg_partial_sum(reg_psum_9_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_0( .activation_in(in_activation_10), .weight_in(reg_weight_9_0), .partial_sum_in(reg_psum_9_0), .reg_activation(reg_activation_10_0), .reg_weight(reg_weight_10_0), .reg_partial_sum(reg_psum_10_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_1( .activation_in(reg_activation_10_0), .weight_in(reg_weight_9_1), .partial_sum_in(reg_psum_9_1), .reg_activation(reg_activation_10_1), .reg_weight(reg_weight_10_1), .reg_partial_sum(reg_psum_10_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_2( .activation_in(reg_activation_10_1), .weight_in(reg_weight_9_2), .partial_sum_in(reg_psum_9_2), .reg_activation(reg_activation_10_2), .reg_weight(reg_weight_10_2), .reg_partial_sum(reg_psum_10_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_3( .activation_in(reg_activation_10_2), .weight_in(reg_weight_9_3), .partial_sum_in(reg_psum_9_3), .reg_activation(reg_activation_10_3), .reg_weight(reg_weight_10_3), .reg_partial_sum(reg_psum_10_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_4( .activation_in(reg_activation_10_3), .weight_in(reg_weight_9_4), .partial_sum_in(reg_psum_9_4), .reg_activation(reg_activation_10_4), .reg_weight(reg_weight_10_4), .reg_partial_sum(reg_psum_10_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_5( .activation_in(reg_activation_10_4), .weight_in(reg_weight_9_5), .partial_sum_in(reg_psum_9_5), .reg_activation(reg_activation_10_5), .reg_weight(reg_weight_10_5), .reg_partial_sum(reg_psum_10_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_6( .activation_in(reg_activation_10_5), .weight_in(reg_weight_9_6), .partial_sum_in(reg_psum_9_6), .reg_activation(reg_activation_10_6), .reg_weight(reg_weight_10_6), .reg_partial_sum(reg_psum_10_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_7( .activation_in(reg_activation_10_6), .weight_in(reg_weight_9_7), .partial_sum_in(reg_psum_9_7), .reg_activation(reg_activation_10_7), .reg_weight(reg_weight_10_7), .reg_partial_sum(reg_psum_10_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_8( .activation_in(reg_activation_10_7), .weight_in(reg_weight_9_8), .partial_sum_in(reg_psum_9_8), .reg_activation(reg_activation_10_8), .reg_weight(reg_weight_10_8), .reg_partial_sum(reg_psum_10_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_9( .activation_in(reg_activation_10_8), .weight_in(reg_weight_9_9), .partial_sum_in(reg_psum_9_9), .reg_activation(reg_activation_10_9), .reg_weight(reg_weight_10_9), .reg_partial_sum(reg_psum_10_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_10( .activation_in(reg_activation_10_9), .weight_in(reg_weight_9_10), .partial_sum_in(reg_psum_9_10), .reg_activation(reg_activation_10_10), .reg_weight(reg_weight_10_10), .reg_partial_sum(reg_psum_10_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_11( .activation_in(reg_activation_10_10), .weight_in(reg_weight_9_11), .partial_sum_in(reg_psum_9_11), .reg_activation(reg_activation_10_11), .reg_weight(reg_weight_10_11), .reg_partial_sum(reg_psum_10_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_12( .activation_in(reg_activation_10_11), .weight_in(reg_weight_9_12), .partial_sum_in(reg_psum_9_12), .reg_activation(reg_activation_10_12), .reg_weight(reg_weight_10_12), .reg_partial_sum(reg_psum_10_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_13( .activation_in(reg_activation_10_12), .weight_in(reg_weight_9_13), .partial_sum_in(reg_psum_9_13), .reg_activation(reg_activation_10_13), .reg_weight(reg_weight_10_13), .reg_partial_sum(reg_psum_10_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_14( .activation_in(reg_activation_10_13), .weight_in(reg_weight_9_14), .partial_sum_in(reg_psum_9_14), .reg_activation(reg_activation_10_14), .reg_weight(reg_weight_10_14), .reg_partial_sum(reg_psum_10_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_15( .activation_in(reg_activation_10_14), .weight_in(reg_weight_9_15), .partial_sum_in(reg_psum_9_15), .reg_activation(reg_activation_10_15), .reg_weight(reg_weight_10_15), .reg_partial_sum(reg_psum_10_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_16( .activation_in(reg_activation_10_15), .weight_in(reg_weight_9_16), .partial_sum_in(reg_psum_9_16), .reg_activation(reg_activation_10_16), .reg_weight(reg_weight_10_16), .reg_partial_sum(reg_psum_10_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_17( .activation_in(reg_activation_10_16), .weight_in(reg_weight_9_17), .partial_sum_in(reg_psum_9_17), .reg_activation(reg_activation_10_17), .reg_weight(reg_weight_10_17), .reg_partial_sum(reg_psum_10_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_18( .activation_in(reg_activation_10_17), .weight_in(reg_weight_9_18), .partial_sum_in(reg_psum_9_18), .reg_activation(reg_activation_10_18), .reg_weight(reg_weight_10_18), .reg_partial_sum(reg_psum_10_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_19( .activation_in(reg_activation_10_18), .weight_in(reg_weight_9_19), .partial_sum_in(reg_psum_9_19), .reg_activation(reg_activation_10_19), .reg_weight(reg_weight_10_19), .reg_partial_sum(reg_psum_10_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_20( .activation_in(reg_activation_10_19), .weight_in(reg_weight_9_20), .partial_sum_in(reg_psum_9_20), .reg_activation(reg_activation_10_20), .reg_weight(reg_weight_10_20), .reg_partial_sum(reg_psum_10_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_21( .activation_in(reg_activation_10_20), .weight_in(reg_weight_9_21), .partial_sum_in(reg_psum_9_21), .reg_activation(reg_activation_10_21), .reg_weight(reg_weight_10_21), .reg_partial_sum(reg_psum_10_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_22( .activation_in(reg_activation_10_21), .weight_in(reg_weight_9_22), .partial_sum_in(reg_psum_9_22), .reg_activation(reg_activation_10_22), .reg_weight(reg_weight_10_22), .reg_partial_sum(reg_psum_10_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_23( .activation_in(reg_activation_10_22), .weight_in(reg_weight_9_23), .partial_sum_in(reg_psum_9_23), .reg_activation(reg_activation_10_23), .reg_weight(reg_weight_10_23), .reg_partial_sum(reg_psum_10_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_24( .activation_in(reg_activation_10_23), .weight_in(reg_weight_9_24), .partial_sum_in(reg_psum_9_24), .reg_activation(reg_activation_10_24), .reg_weight(reg_weight_10_24), .reg_partial_sum(reg_psum_10_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_25( .activation_in(reg_activation_10_24), .weight_in(reg_weight_9_25), .partial_sum_in(reg_psum_9_25), .reg_activation(reg_activation_10_25), .reg_weight(reg_weight_10_25), .reg_partial_sum(reg_psum_10_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_26( .activation_in(reg_activation_10_25), .weight_in(reg_weight_9_26), .partial_sum_in(reg_psum_9_26), .reg_activation(reg_activation_10_26), .reg_weight(reg_weight_10_26), .reg_partial_sum(reg_psum_10_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_27( .activation_in(reg_activation_10_26), .weight_in(reg_weight_9_27), .partial_sum_in(reg_psum_9_27), .reg_activation(reg_activation_10_27), .reg_weight(reg_weight_10_27), .reg_partial_sum(reg_psum_10_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_28( .activation_in(reg_activation_10_27), .weight_in(reg_weight_9_28), .partial_sum_in(reg_psum_9_28), .reg_activation(reg_activation_10_28), .reg_weight(reg_weight_10_28), .reg_partial_sum(reg_psum_10_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_29( .activation_in(reg_activation_10_28), .weight_in(reg_weight_9_29), .partial_sum_in(reg_psum_9_29), .reg_activation(reg_activation_10_29), .reg_weight(reg_weight_10_29), .reg_partial_sum(reg_psum_10_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_30( .activation_in(reg_activation_10_29), .weight_in(reg_weight_9_30), .partial_sum_in(reg_psum_9_30), .reg_activation(reg_activation_10_30), .reg_weight(reg_weight_10_30), .reg_partial_sum(reg_psum_10_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_31( .activation_in(reg_activation_10_30), .weight_in(reg_weight_9_31), .partial_sum_in(reg_psum_9_31), .reg_activation(reg_activation_10_31), .reg_weight(reg_weight_10_31), .reg_partial_sum(reg_psum_10_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_32( .activation_in(reg_activation_10_31), .weight_in(reg_weight_9_32), .partial_sum_in(reg_psum_9_32), .reg_activation(reg_activation_10_32), .reg_weight(reg_weight_10_32), .reg_partial_sum(reg_psum_10_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_33( .activation_in(reg_activation_10_32), .weight_in(reg_weight_9_33), .partial_sum_in(reg_psum_9_33), .reg_activation(reg_activation_10_33), .reg_weight(reg_weight_10_33), .reg_partial_sum(reg_psum_10_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_34( .activation_in(reg_activation_10_33), .weight_in(reg_weight_9_34), .partial_sum_in(reg_psum_9_34), .reg_activation(reg_activation_10_34), .reg_weight(reg_weight_10_34), .reg_partial_sum(reg_psum_10_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_35( .activation_in(reg_activation_10_34), .weight_in(reg_weight_9_35), .partial_sum_in(reg_psum_9_35), .reg_activation(reg_activation_10_35), .reg_weight(reg_weight_10_35), .reg_partial_sum(reg_psum_10_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_36( .activation_in(reg_activation_10_35), .weight_in(reg_weight_9_36), .partial_sum_in(reg_psum_9_36), .reg_activation(reg_activation_10_36), .reg_weight(reg_weight_10_36), .reg_partial_sum(reg_psum_10_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_37( .activation_in(reg_activation_10_36), .weight_in(reg_weight_9_37), .partial_sum_in(reg_psum_9_37), .reg_activation(reg_activation_10_37), .reg_weight(reg_weight_10_37), .reg_partial_sum(reg_psum_10_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_38( .activation_in(reg_activation_10_37), .weight_in(reg_weight_9_38), .partial_sum_in(reg_psum_9_38), .reg_activation(reg_activation_10_38), .reg_weight(reg_weight_10_38), .reg_partial_sum(reg_psum_10_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_39( .activation_in(reg_activation_10_38), .weight_in(reg_weight_9_39), .partial_sum_in(reg_psum_9_39), .reg_activation(reg_activation_10_39), .reg_weight(reg_weight_10_39), .reg_partial_sum(reg_psum_10_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_40( .activation_in(reg_activation_10_39), .weight_in(reg_weight_9_40), .partial_sum_in(reg_psum_9_40), .reg_activation(reg_activation_10_40), .reg_weight(reg_weight_10_40), .reg_partial_sum(reg_psum_10_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_41( .activation_in(reg_activation_10_40), .weight_in(reg_weight_9_41), .partial_sum_in(reg_psum_9_41), .reg_activation(reg_activation_10_41), .reg_weight(reg_weight_10_41), .reg_partial_sum(reg_psum_10_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_42( .activation_in(reg_activation_10_41), .weight_in(reg_weight_9_42), .partial_sum_in(reg_psum_9_42), .reg_activation(reg_activation_10_42), .reg_weight(reg_weight_10_42), .reg_partial_sum(reg_psum_10_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_43( .activation_in(reg_activation_10_42), .weight_in(reg_weight_9_43), .partial_sum_in(reg_psum_9_43), .reg_activation(reg_activation_10_43), .reg_weight(reg_weight_10_43), .reg_partial_sum(reg_psum_10_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_44( .activation_in(reg_activation_10_43), .weight_in(reg_weight_9_44), .partial_sum_in(reg_psum_9_44), .reg_activation(reg_activation_10_44), .reg_weight(reg_weight_10_44), .reg_partial_sum(reg_psum_10_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_45( .activation_in(reg_activation_10_44), .weight_in(reg_weight_9_45), .partial_sum_in(reg_psum_9_45), .reg_activation(reg_activation_10_45), .reg_weight(reg_weight_10_45), .reg_partial_sum(reg_psum_10_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_46( .activation_in(reg_activation_10_45), .weight_in(reg_weight_9_46), .partial_sum_in(reg_psum_9_46), .reg_activation(reg_activation_10_46), .reg_weight(reg_weight_10_46), .reg_partial_sum(reg_psum_10_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_47( .activation_in(reg_activation_10_46), .weight_in(reg_weight_9_47), .partial_sum_in(reg_psum_9_47), .reg_activation(reg_activation_10_47), .reg_weight(reg_weight_10_47), .reg_partial_sum(reg_psum_10_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_48( .activation_in(reg_activation_10_47), .weight_in(reg_weight_9_48), .partial_sum_in(reg_psum_9_48), .reg_activation(reg_activation_10_48), .reg_weight(reg_weight_10_48), .reg_partial_sum(reg_psum_10_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_49( .activation_in(reg_activation_10_48), .weight_in(reg_weight_9_49), .partial_sum_in(reg_psum_9_49), .reg_activation(reg_activation_10_49), .reg_weight(reg_weight_10_49), .reg_partial_sum(reg_psum_10_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_50( .activation_in(reg_activation_10_49), .weight_in(reg_weight_9_50), .partial_sum_in(reg_psum_9_50), .reg_activation(reg_activation_10_50), .reg_weight(reg_weight_10_50), .reg_partial_sum(reg_psum_10_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_51( .activation_in(reg_activation_10_50), .weight_in(reg_weight_9_51), .partial_sum_in(reg_psum_9_51), .reg_activation(reg_activation_10_51), .reg_weight(reg_weight_10_51), .reg_partial_sum(reg_psum_10_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_52( .activation_in(reg_activation_10_51), .weight_in(reg_weight_9_52), .partial_sum_in(reg_psum_9_52), .reg_activation(reg_activation_10_52), .reg_weight(reg_weight_10_52), .reg_partial_sum(reg_psum_10_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_53( .activation_in(reg_activation_10_52), .weight_in(reg_weight_9_53), .partial_sum_in(reg_psum_9_53), .reg_activation(reg_activation_10_53), .reg_weight(reg_weight_10_53), .reg_partial_sum(reg_psum_10_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_54( .activation_in(reg_activation_10_53), .weight_in(reg_weight_9_54), .partial_sum_in(reg_psum_9_54), .reg_activation(reg_activation_10_54), .reg_weight(reg_weight_10_54), .reg_partial_sum(reg_psum_10_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_55( .activation_in(reg_activation_10_54), .weight_in(reg_weight_9_55), .partial_sum_in(reg_psum_9_55), .reg_activation(reg_activation_10_55), .reg_weight(reg_weight_10_55), .reg_partial_sum(reg_psum_10_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_56( .activation_in(reg_activation_10_55), .weight_in(reg_weight_9_56), .partial_sum_in(reg_psum_9_56), .reg_activation(reg_activation_10_56), .reg_weight(reg_weight_10_56), .reg_partial_sum(reg_psum_10_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_57( .activation_in(reg_activation_10_56), .weight_in(reg_weight_9_57), .partial_sum_in(reg_psum_9_57), .reg_activation(reg_activation_10_57), .reg_weight(reg_weight_10_57), .reg_partial_sum(reg_psum_10_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_58( .activation_in(reg_activation_10_57), .weight_in(reg_weight_9_58), .partial_sum_in(reg_psum_9_58), .reg_activation(reg_activation_10_58), .reg_weight(reg_weight_10_58), .reg_partial_sum(reg_psum_10_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_59( .activation_in(reg_activation_10_58), .weight_in(reg_weight_9_59), .partial_sum_in(reg_psum_9_59), .reg_activation(reg_activation_10_59), .reg_weight(reg_weight_10_59), .reg_partial_sum(reg_psum_10_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_60( .activation_in(reg_activation_10_59), .weight_in(reg_weight_9_60), .partial_sum_in(reg_psum_9_60), .reg_activation(reg_activation_10_60), .reg_weight(reg_weight_10_60), .reg_partial_sum(reg_psum_10_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_61( .activation_in(reg_activation_10_60), .weight_in(reg_weight_9_61), .partial_sum_in(reg_psum_9_61), .reg_activation(reg_activation_10_61), .reg_weight(reg_weight_10_61), .reg_partial_sum(reg_psum_10_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_62( .activation_in(reg_activation_10_61), .weight_in(reg_weight_9_62), .partial_sum_in(reg_psum_9_62), .reg_activation(reg_activation_10_62), .reg_weight(reg_weight_10_62), .reg_partial_sum(reg_psum_10_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_63( .activation_in(reg_activation_10_62), .weight_in(reg_weight_9_63), .partial_sum_in(reg_psum_9_63), .reg_weight(reg_weight_10_63), .reg_partial_sum(reg_psum_10_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_0( .activation_in(in_activation_11), .weight_in(reg_weight_10_0), .partial_sum_in(reg_psum_10_0), .reg_activation(reg_activation_11_0), .reg_weight(reg_weight_11_0), .reg_partial_sum(reg_psum_11_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_1( .activation_in(reg_activation_11_0), .weight_in(reg_weight_10_1), .partial_sum_in(reg_psum_10_1), .reg_activation(reg_activation_11_1), .reg_weight(reg_weight_11_1), .reg_partial_sum(reg_psum_11_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_2( .activation_in(reg_activation_11_1), .weight_in(reg_weight_10_2), .partial_sum_in(reg_psum_10_2), .reg_activation(reg_activation_11_2), .reg_weight(reg_weight_11_2), .reg_partial_sum(reg_psum_11_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_3( .activation_in(reg_activation_11_2), .weight_in(reg_weight_10_3), .partial_sum_in(reg_psum_10_3), .reg_activation(reg_activation_11_3), .reg_weight(reg_weight_11_3), .reg_partial_sum(reg_psum_11_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_4( .activation_in(reg_activation_11_3), .weight_in(reg_weight_10_4), .partial_sum_in(reg_psum_10_4), .reg_activation(reg_activation_11_4), .reg_weight(reg_weight_11_4), .reg_partial_sum(reg_psum_11_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_5( .activation_in(reg_activation_11_4), .weight_in(reg_weight_10_5), .partial_sum_in(reg_psum_10_5), .reg_activation(reg_activation_11_5), .reg_weight(reg_weight_11_5), .reg_partial_sum(reg_psum_11_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_6( .activation_in(reg_activation_11_5), .weight_in(reg_weight_10_6), .partial_sum_in(reg_psum_10_6), .reg_activation(reg_activation_11_6), .reg_weight(reg_weight_11_6), .reg_partial_sum(reg_psum_11_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_7( .activation_in(reg_activation_11_6), .weight_in(reg_weight_10_7), .partial_sum_in(reg_psum_10_7), .reg_activation(reg_activation_11_7), .reg_weight(reg_weight_11_7), .reg_partial_sum(reg_psum_11_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_8( .activation_in(reg_activation_11_7), .weight_in(reg_weight_10_8), .partial_sum_in(reg_psum_10_8), .reg_activation(reg_activation_11_8), .reg_weight(reg_weight_11_8), .reg_partial_sum(reg_psum_11_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_9( .activation_in(reg_activation_11_8), .weight_in(reg_weight_10_9), .partial_sum_in(reg_psum_10_9), .reg_activation(reg_activation_11_9), .reg_weight(reg_weight_11_9), .reg_partial_sum(reg_psum_11_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_10( .activation_in(reg_activation_11_9), .weight_in(reg_weight_10_10), .partial_sum_in(reg_psum_10_10), .reg_activation(reg_activation_11_10), .reg_weight(reg_weight_11_10), .reg_partial_sum(reg_psum_11_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_11( .activation_in(reg_activation_11_10), .weight_in(reg_weight_10_11), .partial_sum_in(reg_psum_10_11), .reg_activation(reg_activation_11_11), .reg_weight(reg_weight_11_11), .reg_partial_sum(reg_psum_11_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_12( .activation_in(reg_activation_11_11), .weight_in(reg_weight_10_12), .partial_sum_in(reg_psum_10_12), .reg_activation(reg_activation_11_12), .reg_weight(reg_weight_11_12), .reg_partial_sum(reg_psum_11_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_13( .activation_in(reg_activation_11_12), .weight_in(reg_weight_10_13), .partial_sum_in(reg_psum_10_13), .reg_activation(reg_activation_11_13), .reg_weight(reg_weight_11_13), .reg_partial_sum(reg_psum_11_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_14( .activation_in(reg_activation_11_13), .weight_in(reg_weight_10_14), .partial_sum_in(reg_psum_10_14), .reg_activation(reg_activation_11_14), .reg_weight(reg_weight_11_14), .reg_partial_sum(reg_psum_11_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_15( .activation_in(reg_activation_11_14), .weight_in(reg_weight_10_15), .partial_sum_in(reg_psum_10_15), .reg_activation(reg_activation_11_15), .reg_weight(reg_weight_11_15), .reg_partial_sum(reg_psum_11_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_16( .activation_in(reg_activation_11_15), .weight_in(reg_weight_10_16), .partial_sum_in(reg_psum_10_16), .reg_activation(reg_activation_11_16), .reg_weight(reg_weight_11_16), .reg_partial_sum(reg_psum_11_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_17( .activation_in(reg_activation_11_16), .weight_in(reg_weight_10_17), .partial_sum_in(reg_psum_10_17), .reg_activation(reg_activation_11_17), .reg_weight(reg_weight_11_17), .reg_partial_sum(reg_psum_11_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_18( .activation_in(reg_activation_11_17), .weight_in(reg_weight_10_18), .partial_sum_in(reg_psum_10_18), .reg_activation(reg_activation_11_18), .reg_weight(reg_weight_11_18), .reg_partial_sum(reg_psum_11_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_19( .activation_in(reg_activation_11_18), .weight_in(reg_weight_10_19), .partial_sum_in(reg_psum_10_19), .reg_activation(reg_activation_11_19), .reg_weight(reg_weight_11_19), .reg_partial_sum(reg_psum_11_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_20( .activation_in(reg_activation_11_19), .weight_in(reg_weight_10_20), .partial_sum_in(reg_psum_10_20), .reg_activation(reg_activation_11_20), .reg_weight(reg_weight_11_20), .reg_partial_sum(reg_psum_11_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_21( .activation_in(reg_activation_11_20), .weight_in(reg_weight_10_21), .partial_sum_in(reg_psum_10_21), .reg_activation(reg_activation_11_21), .reg_weight(reg_weight_11_21), .reg_partial_sum(reg_psum_11_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_22( .activation_in(reg_activation_11_21), .weight_in(reg_weight_10_22), .partial_sum_in(reg_psum_10_22), .reg_activation(reg_activation_11_22), .reg_weight(reg_weight_11_22), .reg_partial_sum(reg_psum_11_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_23( .activation_in(reg_activation_11_22), .weight_in(reg_weight_10_23), .partial_sum_in(reg_psum_10_23), .reg_activation(reg_activation_11_23), .reg_weight(reg_weight_11_23), .reg_partial_sum(reg_psum_11_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_24( .activation_in(reg_activation_11_23), .weight_in(reg_weight_10_24), .partial_sum_in(reg_psum_10_24), .reg_activation(reg_activation_11_24), .reg_weight(reg_weight_11_24), .reg_partial_sum(reg_psum_11_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_25( .activation_in(reg_activation_11_24), .weight_in(reg_weight_10_25), .partial_sum_in(reg_psum_10_25), .reg_activation(reg_activation_11_25), .reg_weight(reg_weight_11_25), .reg_partial_sum(reg_psum_11_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_26( .activation_in(reg_activation_11_25), .weight_in(reg_weight_10_26), .partial_sum_in(reg_psum_10_26), .reg_activation(reg_activation_11_26), .reg_weight(reg_weight_11_26), .reg_partial_sum(reg_psum_11_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_27( .activation_in(reg_activation_11_26), .weight_in(reg_weight_10_27), .partial_sum_in(reg_psum_10_27), .reg_activation(reg_activation_11_27), .reg_weight(reg_weight_11_27), .reg_partial_sum(reg_psum_11_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_28( .activation_in(reg_activation_11_27), .weight_in(reg_weight_10_28), .partial_sum_in(reg_psum_10_28), .reg_activation(reg_activation_11_28), .reg_weight(reg_weight_11_28), .reg_partial_sum(reg_psum_11_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_29( .activation_in(reg_activation_11_28), .weight_in(reg_weight_10_29), .partial_sum_in(reg_psum_10_29), .reg_activation(reg_activation_11_29), .reg_weight(reg_weight_11_29), .reg_partial_sum(reg_psum_11_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_30( .activation_in(reg_activation_11_29), .weight_in(reg_weight_10_30), .partial_sum_in(reg_psum_10_30), .reg_activation(reg_activation_11_30), .reg_weight(reg_weight_11_30), .reg_partial_sum(reg_psum_11_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_31( .activation_in(reg_activation_11_30), .weight_in(reg_weight_10_31), .partial_sum_in(reg_psum_10_31), .reg_activation(reg_activation_11_31), .reg_weight(reg_weight_11_31), .reg_partial_sum(reg_psum_11_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_32( .activation_in(reg_activation_11_31), .weight_in(reg_weight_10_32), .partial_sum_in(reg_psum_10_32), .reg_activation(reg_activation_11_32), .reg_weight(reg_weight_11_32), .reg_partial_sum(reg_psum_11_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_33( .activation_in(reg_activation_11_32), .weight_in(reg_weight_10_33), .partial_sum_in(reg_psum_10_33), .reg_activation(reg_activation_11_33), .reg_weight(reg_weight_11_33), .reg_partial_sum(reg_psum_11_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_34( .activation_in(reg_activation_11_33), .weight_in(reg_weight_10_34), .partial_sum_in(reg_psum_10_34), .reg_activation(reg_activation_11_34), .reg_weight(reg_weight_11_34), .reg_partial_sum(reg_psum_11_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_35( .activation_in(reg_activation_11_34), .weight_in(reg_weight_10_35), .partial_sum_in(reg_psum_10_35), .reg_activation(reg_activation_11_35), .reg_weight(reg_weight_11_35), .reg_partial_sum(reg_psum_11_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_36( .activation_in(reg_activation_11_35), .weight_in(reg_weight_10_36), .partial_sum_in(reg_psum_10_36), .reg_activation(reg_activation_11_36), .reg_weight(reg_weight_11_36), .reg_partial_sum(reg_psum_11_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_37( .activation_in(reg_activation_11_36), .weight_in(reg_weight_10_37), .partial_sum_in(reg_psum_10_37), .reg_activation(reg_activation_11_37), .reg_weight(reg_weight_11_37), .reg_partial_sum(reg_psum_11_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_38( .activation_in(reg_activation_11_37), .weight_in(reg_weight_10_38), .partial_sum_in(reg_psum_10_38), .reg_activation(reg_activation_11_38), .reg_weight(reg_weight_11_38), .reg_partial_sum(reg_psum_11_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_39( .activation_in(reg_activation_11_38), .weight_in(reg_weight_10_39), .partial_sum_in(reg_psum_10_39), .reg_activation(reg_activation_11_39), .reg_weight(reg_weight_11_39), .reg_partial_sum(reg_psum_11_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_40( .activation_in(reg_activation_11_39), .weight_in(reg_weight_10_40), .partial_sum_in(reg_psum_10_40), .reg_activation(reg_activation_11_40), .reg_weight(reg_weight_11_40), .reg_partial_sum(reg_psum_11_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_41( .activation_in(reg_activation_11_40), .weight_in(reg_weight_10_41), .partial_sum_in(reg_psum_10_41), .reg_activation(reg_activation_11_41), .reg_weight(reg_weight_11_41), .reg_partial_sum(reg_psum_11_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_42( .activation_in(reg_activation_11_41), .weight_in(reg_weight_10_42), .partial_sum_in(reg_psum_10_42), .reg_activation(reg_activation_11_42), .reg_weight(reg_weight_11_42), .reg_partial_sum(reg_psum_11_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_43( .activation_in(reg_activation_11_42), .weight_in(reg_weight_10_43), .partial_sum_in(reg_psum_10_43), .reg_activation(reg_activation_11_43), .reg_weight(reg_weight_11_43), .reg_partial_sum(reg_psum_11_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_44( .activation_in(reg_activation_11_43), .weight_in(reg_weight_10_44), .partial_sum_in(reg_psum_10_44), .reg_activation(reg_activation_11_44), .reg_weight(reg_weight_11_44), .reg_partial_sum(reg_psum_11_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_45( .activation_in(reg_activation_11_44), .weight_in(reg_weight_10_45), .partial_sum_in(reg_psum_10_45), .reg_activation(reg_activation_11_45), .reg_weight(reg_weight_11_45), .reg_partial_sum(reg_psum_11_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_46( .activation_in(reg_activation_11_45), .weight_in(reg_weight_10_46), .partial_sum_in(reg_psum_10_46), .reg_activation(reg_activation_11_46), .reg_weight(reg_weight_11_46), .reg_partial_sum(reg_psum_11_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_47( .activation_in(reg_activation_11_46), .weight_in(reg_weight_10_47), .partial_sum_in(reg_psum_10_47), .reg_activation(reg_activation_11_47), .reg_weight(reg_weight_11_47), .reg_partial_sum(reg_psum_11_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_48( .activation_in(reg_activation_11_47), .weight_in(reg_weight_10_48), .partial_sum_in(reg_psum_10_48), .reg_activation(reg_activation_11_48), .reg_weight(reg_weight_11_48), .reg_partial_sum(reg_psum_11_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_49( .activation_in(reg_activation_11_48), .weight_in(reg_weight_10_49), .partial_sum_in(reg_psum_10_49), .reg_activation(reg_activation_11_49), .reg_weight(reg_weight_11_49), .reg_partial_sum(reg_psum_11_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_50( .activation_in(reg_activation_11_49), .weight_in(reg_weight_10_50), .partial_sum_in(reg_psum_10_50), .reg_activation(reg_activation_11_50), .reg_weight(reg_weight_11_50), .reg_partial_sum(reg_psum_11_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_51( .activation_in(reg_activation_11_50), .weight_in(reg_weight_10_51), .partial_sum_in(reg_psum_10_51), .reg_activation(reg_activation_11_51), .reg_weight(reg_weight_11_51), .reg_partial_sum(reg_psum_11_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_52( .activation_in(reg_activation_11_51), .weight_in(reg_weight_10_52), .partial_sum_in(reg_psum_10_52), .reg_activation(reg_activation_11_52), .reg_weight(reg_weight_11_52), .reg_partial_sum(reg_psum_11_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_53( .activation_in(reg_activation_11_52), .weight_in(reg_weight_10_53), .partial_sum_in(reg_psum_10_53), .reg_activation(reg_activation_11_53), .reg_weight(reg_weight_11_53), .reg_partial_sum(reg_psum_11_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_54( .activation_in(reg_activation_11_53), .weight_in(reg_weight_10_54), .partial_sum_in(reg_psum_10_54), .reg_activation(reg_activation_11_54), .reg_weight(reg_weight_11_54), .reg_partial_sum(reg_psum_11_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_55( .activation_in(reg_activation_11_54), .weight_in(reg_weight_10_55), .partial_sum_in(reg_psum_10_55), .reg_activation(reg_activation_11_55), .reg_weight(reg_weight_11_55), .reg_partial_sum(reg_psum_11_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_56( .activation_in(reg_activation_11_55), .weight_in(reg_weight_10_56), .partial_sum_in(reg_psum_10_56), .reg_activation(reg_activation_11_56), .reg_weight(reg_weight_11_56), .reg_partial_sum(reg_psum_11_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_57( .activation_in(reg_activation_11_56), .weight_in(reg_weight_10_57), .partial_sum_in(reg_psum_10_57), .reg_activation(reg_activation_11_57), .reg_weight(reg_weight_11_57), .reg_partial_sum(reg_psum_11_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_58( .activation_in(reg_activation_11_57), .weight_in(reg_weight_10_58), .partial_sum_in(reg_psum_10_58), .reg_activation(reg_activation_11_58), .reg_weight(reg_weight_11_58), .reg_partial_sum(reg_psum_11_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_59( .activation_in(reg_activation_11_58), .weight_in(reg_weight_10_59), .partial_sum_in(reg_psum_10_59), .reg_activation(reg_activation_11_59), .reg_weight(reg_weight_11_59), .reg_partial_sum(reg_psum_11_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_60( .activation_in(reg_activation_11_59), .weight_in(reg_weight_10_60), .partial_sum_in(reg_psum_10_60), .reg_activation(reg_activation_11_60), .reg_weight(reg_weight_11_60), .reg_partial_sum(reg_psum_11_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_61( .activation_in(reg_activation_11_60), .weight_in(reg_weight_10_61), .partial_sum_in(reg_psum_10_61), .reg_activation(reg_activation_11_61), .reg_weight(reg_weight_11_61), .reg_partial_sum(reg_psum_11_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_62( .activation_in(reg_activation_11_61), .weight_in(reg_weight_10_62), .partial_sum_in(reg_psum_10_62), .reg_activation(reg_activation_11_62), .reg_weight(reg_weight_11_62), .reg_partial_sum(reg_psum_11_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_63( .activation_in(reg_activation_11_62), .weight_in(reg_weight_10_63), .partial_sum_in(reg_psum_10_63), .reg_weight(reg_weight_11_63), .reg_partial_sum(reg_psum_11_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_0( .activation_in(in_activation_12), .weight_in(reg_weight_11_0), .partial_sum_in(reg_psum_11_0), .reg_activation(reg_activation_12_0), .reg_weight(reg_weight_12_0), .reg_partial_sum(reg_psum_12_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_1( .activation_in(reg_activation_12_0), .weight_in(reg_weight_11_1), .partial_sum_in(reg_psum_11_1), .reg_activation(reg_activation_12_1), .reg_weight(reg_weight_12_1), .reg_partial_sum(reg_psum_12_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_2( .activation_in(reg_activation_12_1), .weight_in(reg_weight_11_2), .partial_sum_in(reg_psum_11_2), .reg_activation(reg_activation_12_2), .reg_weight(reg_weight_12_2), .reg_partial_sum(reg_psum_12_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_3( .activation_in(reg_activation_12_2), .weight_in(reg_weight_11_3), .partial_sum_in(reg_psum_11_3), .reg_activation(reg_activation_12_3), .reg_weight(reg_weight_12_3), .reg_partial_sum(reg_psum_12_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_4( .activation_in(reg_activation_12_3), .weight_in(reg_weight_11_4), .partial_sum_in(reg_psum_11_4), .reg_activation(reg_activation_12_4), .reg_weight(reg_weight_12_4), .reg_partial_sum(reg_psum_12_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_5( .activation_in(reg_activation_12_4), .weight_in(reg_weight_11_5), .partial_sum_in(reg_psum_11_5), .reg_activation(reg_activation_12_5), .reg_weight(reg_weight_12_5), .reg_partial_sum(reg_psum_12_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_6( .activation_in(reg_activation_12_5), .weight_in(reg_weight_11_6), .partial_sum_in(reg_psum_11_6), .reg_activation(reg_activation_12_6), .reg_weight(reg_weight_12_6), .reg_partial_sum(reg_psum_12_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_7( .activation_in(reg_activation_12_6), .weight_in(reg_weight_11_7), .partial_sum_in(reg_psum_11_7), .reg_activation(reg_activation_12_7), .reg_weight(reg_weight_12_7), .reg_partial_sum(reg_psum_12_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_8( .activation_in(reg_activation_12_7), .weight_in(reg_weight_11_8), .partial_sum_in(reg_psum_11_8), .reg_activation(reg_activation_12_8), .reg_weight(reg_weight_12_8), .reg_partial_sum(reg_psum_12_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_9( .activation_in(reg_activation_12_8), .weight_in(reg_weight_11_9), .partial_sum_in(reg_psum_11_9), .reg_activation(reg_activation_12_9), .reg_weight(reg_weight_12_9), .reg_partial_sum(reg_psum_12_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_10( .activation_in(reg_activation_12_9), .weight_in(reg_weight_11_10), .partial_sum_in(reg_psum_11_10), .reg_activation(reg_activation_12_10), .reg_weight(reg_weight_12_10), .reg_partial_sum(reg_psum_12_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_11( .activation_in(reg_activation_12_10), .weight_in(reg_weight_11_11), .partial_sum_in(reg_psum_11_11), .reg_activation(reg_activation_12_11), .reg_weight(reg_weight_12_11), .reg_partial_sum(reg_psum_12_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_12( .activation_in(reg_activation_12_11), .weight_in(reg_weight_11_12), .partial_sum_in(reg_psum_11_12), .reg_activation(reg_activation_12_12), .reg_weight(reg_weight_12_12), .reg_partial_sum(reg_psum_12_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_13( .activation_in(reg_activation_12_12), .weight_in(reg_weight_11_13), .partial_sum_in(reg_psum_11_13), .reg_activation(reg_activation_12_13), .reg_weight(reg_weight_12_13), .reg_partial_sum(reg_psum_12_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_14( .activation_in(reg_activation_12_13), .weight_in(reg_weight_11_14), .partial_sum_in(reg_psum_11_14), .reg_activation(reg_activation_12_14), .reg_weight(reg_weight_12_14), .reg_partial_sum(reg_psum_12_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_15( .activation_in(reg_activation_12_14), .weight_in(reg_weight_11_15), .partial_sum_in(reg_psum_11_15), .reg_activation(reg_activation_12_15), .reg_weight(reg_weight_12_15), .reg_partial_sum(reg_psum_12_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_16( .activation_in(reg_activation_12_15), .weight_in(reg_weight_11_16), .partial_sum_in(reg_psum_11_16), .reg_activation(reg_activation_12_16), .reg_weight(reg_weight_12_16), .reg_partial_sum(reg_psum_12_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_17( .activation_in(reg_activation_12_16), .weight_in(reg_weight_11_17), .partial_sum_in(reg_psum_11_17), .reg_activation(reg_activation_12_17), .reg_weight(reg_weight_12_17), .reg_partial_sum(reg_psum_12_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_18( .activation_in(reg_activation_12_17), .weight_in(reg_weight_11_18), .partial_sum_in(reg_psum_11_18), .reg_activation(reg_activation_12_18), .reg_weight(reg_weight_12_18), .reg_partial_sum(reg_psum_12_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_19( .activation_in(reg_activation_12_18), .weight_in(reg_weight_11_19), .partial_sum_in(reg_psum_11_19), .reg_activation(reg_activation_12_19), .reg_weight(reg_weight_12_19), .reg_partial_sum(reg_psum_12_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_20( .activation_in(reg_activation_12_19), .weight_in(reg_weight_11_20), .partial_sum_in(reg_psum_11_20), .reg_activation(reg_activation_12_20), .reg_weight(reg_weight_12_20), .reg_partial_sum(reg_psum_12_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_21( .activation_in(reg_activation_12_20), .weight_in(reg_weight_11_21), .partial_sum_in(reg_psum_11_21), .reg_activation(reg_activation_12_21), .reg_weight(reg_weight_12_21), .reg_partial_sum(reg_psum_12_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_22( .activation_in(reg_activation_12_21), .weight_in(reg_weight_11_22), .partial_sum_in(reg_psum_11_22), .reg_activation(reg_activation_12_22), .reg_weight(reg_weight_12_22), .reg_partial_sum(reg_psum_12_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_23( .activation_in(reg_activation_12_22), .weight_in(reg_weight_11_23), .partial_sum_in(reg_psum_11_23), .reg_activation(reg_activation_12_23), .reg_weight(reg_weight_12_23), .reg_partial_sum(reg_psum_12_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_24( .activation_in(reg_activation_12_23), .weight_in(reg_weight_11_24), .partial_sum_in(reg_psum_11_24), .reg_activation(reg_activation_12_24), .reg_weight(reg_weight_12_24), .reg_partial_sum(reg_psum_12_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_25( .activation_in(reg_activation_12_24), .weight_in(reg_weight_11_25), .partial_sum_in(reg_psum_11_25), .reg_activation(reg_activation_12_25), .reg_weight(reg_weight_12_25), .reg_partial_sum(reg_psum_12_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_26( .activation_in(reg_activation_12_25), .weight_in(reg_weight_11_26), .partial_sum_in(reg_psum_11_26), .reg_activation(reg_activation_12_26), .reg_weight(reg_weight_12_26), .reg_partial_sum(reg_psum_12_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_27( .activation_in(reg_activation_12_26), .weight_in(reg_weight_11_27), .partial_sum_in(reg_psum_11_27), .reg_activation(reg_activation_12_27), .reg_weight(reg_weight_12_27), .reg_partial_sum(reg_psum_12_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_28( .activation_in(reg_activation_12_27), .weight_in(reg_weight_11_28), .partial_sum_in(reg_psum_11_28), .reg_activation(reg_activation_12_28), .reg_weight(reg_weight_12_28), .reg_partial_sum(reg_psum_12_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_29( .activation_in(reg_activation_12_28), .weight_in(reg_weight_11_29), .partial_sum_in(reg_psum_11_29), .reg_activation(reg_activation_12_29), .reg_weight(reg_weight_12_29), .reg_partial_sum(reg_psum_12_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_30( .activation_in(reg_activation_12_29), .weight_in(reg_weight_11_30), .partial_sum_in(reg_psum_11_30), .reg_activation(reg_activation_12_30), .reg_weight(reg_weight_12_30), .reg_partial_sum(reg_psum_12_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_31( .activation_in(reg_activation_12_30), .weight_in(reg_weight_11_31), .partial_sum_in(reg_psum_11_31), .reg_activation(reg_activation_12_31), .reg_weight(reg_weight_12_31), .reg_partial_sum(reg_psum_12_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_32( .activation_in(reg_activation_12_31), .weight_in(reg_weight_11_32), .partial_sum_in(reg_psum_11_32), .reg_activation(reg_activation_12_32), .reg_weight(reg_weight_12_32), .reg_partial_sum(reg_psum_12_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_33( .activation_in(reg_activation_12_32), .weight_in(reg_weight_11_33), .partial_sum_in(reg_psum_11_33), .reg_activation(reg_activation_12_33), .reg_weight(reg_weight_12_33), .reg_partial_sum(reg_psum_12_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_34( .activation_in(reg_activation_12_33), .weight_in(reg_weight_11_34), .partial_sum_in(reg_psum_11_34), .reg_activation(reg_activation_12_34), .reg_weight(reg_weight_12_34), .reg_partial_sum(reg_psum_12_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_35( .activation_in(reg_activation_12_34), .weight_in(reg_weight_11_35), .partial_sum_in(reg_psum_11_35), .reg_activation(reg_activation_12_35), .reg_weight(reg_weight_12_35), .reg_partial_sum(reg_psum_12_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_36( .activation_in(reg_activation_12_35), .weight_in(reg_weight_11_36), .partial_sum_in(reg_psum_11_36), .reg_activation(reg_activation_12_36), .reg_weight(reg_weight_12_36), .reg_partial_sum(reg_psum_12_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_37( .activation_in(reg_activation_12_36), .weight_in(reg_weight_11_37), .partial_sum_in(reg_psum_11_37), .reg_activation(reg_activation_12_37), .reg_weight(reg_weight_12_37), .reg_partial_sum(reg_psum_12_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_38( .activation_in(reg_activation_12_37), .weight_in(reg_weight_11_38), .partial_sum_in(reg_psum_11_38), .reg_activation(reg_activation_12_38), .reg_weight(reg_weight_12_38), .reg_partial_sum(reg_psum_12_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_39( .activation_in(reg_activation_12_38), .weight_in(reg_weight_11_39), .partial_sum_in(reg_psum_11_39), .reg_activation(reg_activation_12_39), .reg_weight(reg_weight_12_39), .reg_partial_sum(reg_psum_12_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_40( .activation_in(reg_activation_12_39), .weight_in(reg_weight_11_40), .partial_sum_in(reg_psum_11_40), .reg_activation(reg_activation_12_40), .reg_weight(reg_weight_12_40), .reg_partial_sum(reg_psum_12_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_41( .activation_in(reg_activation_12_40), .weight_in(reg_weight_11_41), .partial_sum_in(reg_psum_11_41), .reg_activation(reg_activation_12_41), .reg_weight(reg_weight_12_41), .reg_partial_sum(reg_psum_12_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_42( .activation_in(reg_activation_12_41), .weight_in(reg_weight_11_42), .partial_sum_in(reg_psum_11_42), .reg_activation(reg_activation_12_42), .reg_weight(reg_weight_12_42), .reg_partial_sum(reg_psum_12_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_43( .activation_in(reg_activation_12_42), .weight_in(reg_weight_11_43), .partial_sum_in(reg_psum_11_43), .reg_activation(reg_activation_12_43), .reg_weight(reg_weight_12_43), .reg_partial_sum(reg_psum_12_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_44( .activation_in(reg_activation_12_43), .weight_in(reg_weight_11_44), .partial_sum_in(reg_psum_11_44), .reg_activation(reg_activation_12_44), .reg_weight(reg_weight_12_44), .reg_partial_sum(reg_psum_12_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_45( .activation_in(reg_activation_12_44), .weight_in(reg_weight_11_45), .partial_sum_in(reg_psum_11_45), .reg_activation(reg_activation_12_45), .reg_weight(reg_weight_12_45), .reg_partial_sum(reg_psum_12_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_46( .activation_in(reg_activation_12_45), .weight_in(reg_weight_11_46), .partial_sum_in(reg_psum_11_46), .reg_activation(reg_activation_12_46), .reg_weight(reg_weight_12_46), .reg_partial_sum(reg_psum_12_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_47( .activation_in(reg_activation_12_46), .weight_in(reg_weight_11_47), .partial_sum_in(reg_psum_11_47), .reg_activation(reg_activation_12_47), .reg_weight(reg_weight_12_47), .reg_partial_sum(reg_psum_12_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_48( .activation_in(reg_activation_12_47), .weight_in(reg_weight_11_48), .partial_sum_in(reg_psum_11_48), .reg_activation(reg_activation_12_48), .reg_weight(reg_weight_12_48), .reg_partial_sum(reg_psum_12_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_49( .activation_in(reg_activation_12_48), .weight_in(reg_weight_11_49), .partial_sum_in(reg_psum_11_49), .reg_activation(reg_activation_12_49), .reg_weight(reg_weight_12_49), .reg_partial_sum(reg_psum_12_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_50( .activation_in(reg_activation_12_49), .weight_in(reg_weight_11_50), .partial_sum_in(reg_psum_11_50), .reg_activation(reg_activation_12_50), .reg_weight(reg_weight_12_50), .reg_partial_sum(reg_psum_12_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_51( .activation_in(reg_activation_12_50), .weight_in(reg_weight_11_51), .partial_sum_in(reg_psum_11_51), .reg_activation(reg_activation_12_51), .reg_weight(reg_weight_12_51), .reg_partial_sum(reg_psum_12_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_52( .activation_in(reg_activation_12_51), .weight_in(reg_weight_11_52), .partial_sum_in(reg_psum_11_52), .reg_activation(reg_activation_12_52), .reg_weight(reg_weight_12_52), .reg_partial_sum(reg_psum_12_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_53( .activation_in(reg_activation_12_52), .weight_in(reg_weight_11_53), .partial_sum_in(reg_psum_11_53), .reg_activation(reg_activation_12_53), .reg_weight(reg_weight_12_53), .reg_partial_sum(reg_psum_12_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_54( .activation_in(reg_activation_12_53), .weight_in(reg_weight_11_54), .partial_sum_in(reg_psum_11_54), .reg_activation(reg_activation_12_54), .reg_weight(reg_weight_12_54), .reg_partial_sum(reg_psum_12_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_55( .activation_in(reg_activation_12_54), .weight_in(reg_weight_11_55), .partial_sum_in(reg_psum_11_55), .reg_activation(reg_activation_12_55), .reg_weight(reg_weight_12_55), .reg_partial_sum(reg_psum_12_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_56( .activation_in(reg_activation_12_55), .weight_in(reg_weight_11_56), .partial_sum_in(reg_psum_11_56), .reg_activation(reg_activation_12_56), .reg_weight(reg_weight_12_56), .reg_partial_sum(reg_psum_12_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_57( .activation_in(reg_activation_12_56), .weight_in(reg_weight_11_57), .partial_sum_in(reg_psum_11_57), .reg_activation(reg_activation_12_57), .reg_weight(reg_weight_12_57), .reg_partial_sum(reg_psum_12_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_58( .activation_in(reg_activation_12_57), .weight_in(reg_weight_11_58), .partial_sum_in(reg_psum_11_58), .reg_activation(reg_activation_12_58), .reg_weight(reg_weight_12_58), .reg_partial_sum(reg_psum_12_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_59( .activation_in(reg_activation_12_58), .weight_in(reg_weight_11_59), .partial_sum_in(reg_psum_11_59), .reg_activation(reg_activation_12_59), .reg_weight(reg_weight_12_59), .reg_partial_sum(reg_psum_12_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_60( .activation_in(reg_activation_12_59), .weight_in(reg_weight_11_60), .partial_sum_in(reg_psum_11_60), .reg_activation(reg_activation_12_60), .reg_weight(reg_weight_12_60), .reg_partial_sum(reg_psum_12_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_61( .activation_in(reg_activation_12_60), .weight_in(reg_weight_11_61), .partial_sum_in(reg_psum_11_61), .reg_activation(reg_activation_12_61), .reg_weight(reg_weight_12_61), .reg_partial_sum(reg_psum_12_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_62( .activation_in(reg_activation_12_61), .weight_in(reg_weight_11_62), .partial_sum_in(reg_psum_11_62), .reg_activation(reg_activation_12_62), .reg_weight(reg_weight_12_62), .reg_partial_sum(reg_psum_12_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_63( .activation_in(reg_activation_12_62), .weight_in(reg_weight_11_63), .partial_sum_in(reg_psum_11_63), .reg_weight(reg_weight_12_63), .reg_partial_sum(reg_psum_12_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_0( .activation_in(in_activation_13), .weight_in(reg_weight_12_0), .partial_sum_in(reg_psum_12_0), .reg_activation(reg_activation_13_0), .reg_weight(reg_weight_13_0), .reg_partial_sum(reg_psum_13_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_1( .activation_in(reg_activation_13_0), .weight_in(reg_weight_12_1), .partial_sum_in(reg_psum_12_1), .reg_activation(reg_activation_13_1), .reg_weight(reg_weight_13_1), .reg_partial_sum(reg_psum_13_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_2( .activation_in(reg_activation_13_1), .weight_in(reg_weight_12_2), .partial_sum_in(reg_psum_12_2), .reg_activation(reg_activation_13_2), .reg_weight(reg_weight_13_2), .reg_partial_sum(reg_psum_13_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_3( .activation_in(reg_activation_13_2), .weight_in(reg_weight_12_3), .partial_sum_in(reg_psum_12_3), .reg_activation(reg_activation_13_3), .reg_weight(reg_weight_13_3), .reg_partial_sum(reg_psum_13_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_4( .activation_in(reg_activation_13_3), .weight_in(reg_weight_12_4), .partial_sum_in(reg_psum_12_4), .reg_activation(reg_activation_13_4), .reg_weight(reg_weight_13_4), .reg_partial_sum(reg_psum_13_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_5( .activation_in(reg_activation_13_4), .weight_in(reg_weight_12_5), .partial_sum_in(reg_psum_12_5), .reg_activation(reg_activation_13_5), .reg_weight(reg_weight_13_5), .reg_partial_sum(reg_psum_13_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_6( .activation_in(reg_activation_13_5), .weight_in(reg_weight_12_6), .partial_sum_in(reg_psum_12_6), .reg_activation(reg_activation_13_6), .reg_weight(reg_weight_13_6), .reg_partial_sum(reg_psum_13_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_7( .activation_in(reg_activation_13_6), .weight_in(reg_weight_12_7), .partial_sum_in(reg_psum_12_7), .reg_activation(reg_activation_13_7), .reg_weight(reg_weight_13_7), .reg_partial_sum(reg_psum_13_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_8( .activation_in(reg_activation_13_7), .weight_in(reg_weight_12_8), .partial_sum_in(reg_psum_12_8), .reg_activation(reg_activation_13_8), .reg_weight(reg_weight_13_8), .reg_partial_sum(reg_psum_13_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_9( .activation_in(reg_activation_13_8), .weight_in(reg_weight_12_9), .partial_sum_in(reg_psum_12_9), .reg_activation(reg_activation_13_9), .reg_weight(reg_weight_13_9), .reg_partial_sum(reg_psum_13_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_10( .activation_in(reg_activation_13_9), .weight_in(reg_weight_12_10), .partial_sum_in(reg_psum_12_10), .reg_activation(reg_activation_13_10), .reg_weight(reg_weight_13_10), .reg_partial_sum(reg_psum_13_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_11( .activation_in(reg_activation_13_10), .weight_in(reg_weight_12_11), .partial_sum_in(reg_psum_12_11), .reg_activation(reg_activation_13_11), .reg_weight(reg_weight_13_11), .reg_partial_sum(reg_psum_13_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_12( .activation_in(reg_activation_13_11), .weight_in(reg_weight_12_12), .partial_sum_in(reg_psum_12_12), .reg_activation(reg_activation_13_12), .reg_weight(reg_weight_13_12), .reg_partial_sum(reg_psum_13_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_13( .activation_in(reg_activation_13_12), .weight_in(reg_weight_12_13), .partial_sum_in(reg_psum_12_13), .reg_activation(reg_activation_13_13), .reg_weight(reg_weight_13_13), .reg_partial_sum(reg_psum_13_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_14( .activation_in(reg_activation_13_13), .weight_in(reg_weight_12_14), .partial_sum_in(reg_psum_12_14), .reg_activation(reg_activation_13_14), .reg_weight(reg_weight_13_14), .reg_partial_sum(reg_psum_13_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_15( .activation_in(reg_activation_13_14), .weight_in(reg_weight_12_15), .partial_sum_in(reg_psum_12_15), .reg_activation(reg_activation_13_15), .reg_weight(reg_weight_13_15), .reg_partial_sum(reg_psum_13_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_16( .activation_in(reg_activation_13_15), .weight_in(reg_weight_12_16), .partial_sum_in(reg_psum_12_16), .reg_activation(reg_activation_13_16), .reg_weight(reg_weight_13_16), .reg_partial_sum(reg_psum_13_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_17( .activation_in(reg_activation_13_16), .weight_in(reg_weight_12_17), .partial_sum_in(reg_psum_12_17), .reg_activation(reg_activation_13_17), .reg_weight(reg_weight_13_17), .reg_partial_sum(reg_psum_13_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_18( .activation_in(reg_activation_13_17), .weight_in(reg_weight_12_18), .partial_sum_in(reg_psum_12_18), .reg_activation(reg_activation_13_18), .reg_weight(reg_weight_13_18), .reg_partial_sum(reg_psum_13_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_19( .activation_in(reg_activation_13_18), .weight_in(reg_weight_12_19), .partial_sum_in(reg_psum_12_19), .reg_activation(reg_activation_13_19), .reg_weight(reg_weight_13_19), .reg_partial_sum(reg_psum_13_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_20( .activation_in(reg_activation_13_19), .weight_in(reg_weight_12_20), .partial_sum_in(reg_psum_12_20), .reg_activation(reg_activation_13_20), .reg_weight(reg_weight_13_20), .reg_partial_sum(reg_psum_13_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_21( .activation_in(reg_activation_13_20), .weight_in(reg_weight_12_21), .partial_sum_in(reg_psum_12_21), .reg_activation(reg_activation_13_21), .reg_weight(reg_weight_13_21), .reg_partial_sum(reg_psum_13_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_22( .activation_in(reg_activation_13_21), .weight_in(reg_weight_12_22), .partial_sum_in(reg_psum_12_22), .reg_activation(reg_activation_13_22), .reg_weight(reg_weight_13_22), .reg_partial_sum(reg_psum_13_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_23( .activation_in(reg_activation_13_22), .weight_in(reg_weight_12_23), .partial_sum_in(reg_psum_12_23), .reg_activation(reg_activation_13_23), .reg_weight(reg_weight_13_23), .reg_partial_sum(reg_psum_13_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_24( .activation_in(reg_activation_13_23), .weight_in(reg_weight_12_24), .partial_sum_in(reg_psum_12_24), .reg_activation(reg_activation_13_24), .reg_weight(reg_weight_13_24), .reg_partial_sum(reg_psum_13_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_25( .activation_in(reg_activation_13_24), .weight_in(reg_weight_12_25), .partial_sum_in(reg_psum_12_25), .reg_activation(reg_activation_13_25), .reg_weight(reg_weight_13_25), .reg_partial_sum(reg_psum_13_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_26( .activation_in(reg_activation_13_25), .weight_in(reg_weight_12_26), .partial_sum_in(reg_psum_12_26), .reg_activation(reg_activation_13_26), .reg_weight(reg_weight_13_26), .reg_partial_sum(reg_psum_13_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_27( .activation_in(reg_activation_13_26), .weight_in(reg_weight_12_27), .partial_sum_in(reg_psum_12_27), .reg_activation(reg_activation_13_27), .reg_weight(reg_weight_13_27), .reg_partial_sum(reg_psum_13_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_28( .activation_in(reg_activation_13_27), .weight_in(reg_weight_12_28), .partial_sum_in(reg_psum_12_28), .reg_activation(reg_activation_13_28), .reg_weight(reg_weight_13_28), .reg_partial_sum(reg_psum_13_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_29( .activation_in(reg_activation_13_28), .weight_in(reg_weight_12_29), .partial_sum_in(reg_psum_12_29), .reg_activation(reg_activation_13_29), .reg_weight(reg_weight_13_29), .reg_partial_sum(reg_psum_13_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_30( .activation_in(reg_activation_13_29), .weight_in(reg_weight_12_30), .partial_sum_in(reg_psum_12_30), .reg_activation(reg_activation_13_30), .reg_weight(reg_weight_13_30), .reg_partial_sum(reg_psum_13_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_31( .activation_in(reg_activation_13_30), .weight_in(reg_weight_12_31), .partial_sum_in(reg_psum_12_31), .reg_activation(reg_activation_13_31), .reg_weight(reg_weight_13_31), .reg_partial_sum(reg_psum_13_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_32( .activation_in(reg_activation_13_31), .weight_in(reg_weight_12_32), .partial_sum_in(reg_psum_12_32), .reg_activation(reg_activation_13_32), .reg_weight(reg_weight_13_32), .reg_partial_sum(reg_psum_13_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_33( .activation_in(reg_activation_13_32), .weight_in(reg_weight_12_33), .partial_sum_in(reg_psum_12_33), .reg_activation(reg_activation_13_33), .reg_weight(reg_weight_13_33), .reg_partial_sum(reg_psum_13_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_34( .activation_in(reg_activation_13_33), .weight_in(reg_weight_12_34), .partial_sum_in(reg_psum_12_34), .reg_activation(reg_activation_13_34), .reg_weight(reg_weight_13_34), .reg_partial_sum(reg_psum_13_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_35( .activation_in(reg_activation_13_34), .weight_in(reg_weight_12_35), .partial_sum_in(reg_psum_12_35), .reg_activation(reg_activation_13_35), .reg_weight(reg_weight_13_35), .reg_partial_sum(reg_psum_13_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_36( .activation_in(reg_activation_13_35), .weight_in(reg_weight_12_36), .partial_sum_in(reg_psum_12_36), .reg_activation(reg_activation_13_36), .reg_weight(reg_weight_13_36), .reg_partial_sum(reg_psum_13_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_37( .activation_in(reg_activation_13_36), .weight_in(reg_weight_12_37), .partial_sum_in(reg_psum_12_37), .reg_activation(reg_activation_13_37), .reg_weight(reg_weight_13_37), .reg_partial_sum(reg_psum_13_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_38( .activation_in(reg_activation_13_37), .weight_in(reg_weight_12_38), .partial_sum_in(reg_psum_12_38), .reg_activation(reg_activation_13_38), .reg_weight(reg_weight_13_38), .reg_partial_sum(reg_psum_13_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_39( .activation_in(reg_activation_13_38), .weight_in(reg_weight_12_39), .partial_sum_in(reg_psum_12_39), .reg_activation(reg_activation_13_39), .reg_weight(reg_weight_13_39), .reg_partial_sum(reg_psum_13_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_40( .activation_in(reg_activation_13_39), .weight_in(reg_weight_12_40), .partial_sum_in(reg_psum_12_40), .reg_activation(reg_activation_13_40), .reg_weight(reg_weight_13_40), .reg_partial_sum(reg_psum_13_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_41( .activation_in(reg_activation_13_40), .weight_in(reg_weight_12_41), .partial_sum_in(reg_psum_12_41), .reg_activation(reg_activation_13_41), .reg_weight(reg_weight_13_41), .reg_partial_sum(reg_psum_13_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_42( .activation_in(reg_activation_13_41), .weight_in(reg_weight_12_42), .partial_sum_in(reg_psum_12_42), .reg_activation(reg_activation_13_42), .reg_weight(reg_weight_13_42), .reg_partial_sum(reg_psum_13_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_43( .activation_in(reg_activation_13_42), .weight_in(reg_weight_12_43), .partial_sum_in(reg_psum_12_43), .reg_activation(reg_activation_13_43), .reg_weight(reg_weight_13_43), .reg_partial_sum(reg_psum_13_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_44( .activation_in(reg_activation_13_43), .weight_in(reg_weight_12_44), .partial_sum_in(reg_psum_12_44), .reg_activation(reg_activation_13_44), .reg_weight(reg_weight_13_44), .reg_partial_sum(reg_psum_13_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_45( .activation_in(reg_activation_13_44), .weight_in(reg_weight_12_45), .partial_sum_in(reg_psum_12_45), .reg_activation(reg_activation_13_45), .reg_weight(reg_weight_13_45), .reg_partial_sum(reg_psum_13_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_46( .activation_in(reg_activation_13_45), .weight_in(reg_weight_12_46), .partial_sum_in(reg_psum_12_46), .reg_activation(reg_activation_13_46), .reg_weight(reg_weight_13_46), .reg_partial_sum(reg_psum_13_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_47( .activation_in(reg_activation_13_46), .weight_in(reg_weight_12_47), .partial_sum_in(reg_psum_12_47), .reg_activation(reg_activation_13_47), .reg_weight(reg_weight_13_47), .reg_partial_sum(reg_psum_13_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_48( .activation_in(reg_activation_13_47), .weight_in(reg_weight_12_48), .partial_sum_in(reg_psum_12_48), .reg_activation(reg_activation_13_48), .reg_weight(reg_weight_13_48), .reg_partial_sum(reg_psum_13_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_49( .activation_in(reg_activation_13_48), .weight_in(reg_weight_12_49), .partial_sum_in(reg_psum_12_49), .reg_activation(reg_activation_13_49), .reg_weight(reg_weight_13_49), .reg_partial_sum(reg_psum_13_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_50( .activation_in(reg_activation_13_49), .weight_in(reg_weight_12_50), .partial_sum_in(reg_psum_12_50), .reg_activation(reg_activation_13_50), .reg_weight(reg_weight_13_50), .reg_partial_sum(reg_psum_13_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_51( .activation_in(reg_activation_13_50), .weight_in(reg_weight_12_51), .partial_sum_in(reg_psum_12_51), .reg_activation(reg_activation_13_51), .reg_weight(reg_weight_13_51), .reg_partial_sum(reg_psum_13_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_52( .activation_in(reg_activation_13_51), .weight_in(reg_weight_12_52), .partial_sum_in(reg_psum_12_52), .reg_activation(reg_activation_13_52), .reg_weight(reg_weight_13_52), .reg_partial_sum(reg_psum_13_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_53( .activation_in(reg_activation_13_52), .weight_in(reg_weight_12_53), .partial_sum_in(reg_psum_12_53), .reg_activation(reg_activation_13_53), .reg_weight(reg_weight_13_53), .reg_partial_sum(reg_psum_13_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_54( .activation_in(reg_activation_13_53), .weight_in(reg_weight_12_54), .partial_sum_in(reg_psum_12_54), .reg_activation(reg_activation_13_54), .reg_weight(reg_weight_13_54), .reg_partial_sum(reg_psum_13_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_55( .activation_in(reg_activation_13_54), .weight_in(reg_weight_12_55), .partial_sum_in(reg_psum_12_55), .reg_activation(reg_activation_13_55), .reg_weight(reg_weight_13_55), .reg_partial_sum(reg_psum_13_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_56( .activation_in(reg_activation_13_55), .weight_in(reg_weight_12_56), .partial_sum_in(reg_psum_12_56), .reg_activation(reg_activation_13_56), .reg_weight(reg_weight_13_56), .reg_partial_sum(reg_psum_13_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_57( .activation_in(reg_activation_13_56), .weight_in(reg_weight_12_57), .partial_sum_in(reg_psum_12_57), .reg_activation(reg_activation_13_57), .reg_weight(reg_weight_13_57), .reg_partial_sum(reg_psum_13_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_58( .activation_in(reg_activation_13_57), .weight_in(reg_weight_12_58), .partial_sum_in(reg_psum_12_58), .reg_activation(reg_activation_13_58), .reg_weight(reg_weight_13_58), .reg_partial_sum(reg_psum_13_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_59( .activation_in(reg_activation_13_58), .weight_in(reg_weight_12_59), .partial_sum_in(reg_psum_12_59), .reg_activation(reg_activation_13_59), .reg_weight(reg_weight_13_59), .reg_partial_sum(reg_psum_13_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_60( .activation_in(reg_activation_13_59), .weight_in(reg_weight_12_60), .partial_sum_in(reg_psum_12_60), .reg_activation(reg_activation_13_60), .reg_weight(reg_weight_13_60), .reg_partial_sum(reg_psum_13_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_61( .activation_in(reg_activation_13_60), .weight_in(reg_weight_12_61), .partial_sum_in(reg_psum_12_61), .reg_activation(reg_activation_13_61), .reg_weight(reg_weight_13_61), .reg_partial_sum(reg_psum_13_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_62( .activation_in(reg_activation_13_61), .weight_in(reg_weight_12_62), .partial_sum_in(reg_psum_12_62), .reg_activation(reg_activation_13_62), .reg_weight(reg_weight_13_62), .reg_partial_sum(reg_psum_13_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_63( .activation_in(reg_activation_13_62), .weight_in(reg_weight_12_63), .partial_sum_in(reg_psum_12_63), .reg_weight(reg_weight_13_63), .reg_partial_sum(reg_psum_13_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_0( .activation_in(in_activation_14), .weight_in(reg_weight_13_0), .partial_sum_in(reg_psum_13_0), .reg_activation(reg_activation_14_0), .reg_weight(reg_weight_14_0), .reg_partial_sum(reg_psum_14_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_1( .activation_in(reg_activation_14_0), .weight_in(reg_weight_13_1), .partial_sum_in(reg_psum_13_1), .reg_activation(reg_activation_14_1), .reg_weight(reg_weight_14_1), .reg_partial_sum(reg_psum_14_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_2( .activation_in(reg_activation_14_1), .weight_in(reg_weight_13_2), .partial_sum_in(reg_psum_13_2), .reg_activation(reg_activation_14_2), .reg_weight(reg_weight_14_2), .reg_partial_sum(reg_psum_14_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_3( .activation_in(reg_activation_14_2), .weight_in(reg_weight_13_3), .partial_sum_in(reg_psum_13_3), .reg_activation(reg_activation_14_3), .reg_weight(reg_weight_14_3), .reg_partial_sum(reg_psum_14_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_4( .activation_in(reg_activation_14_3), .weight_in(reg_weight_13_4), .partial_sum_in(reg_psum_13_4), .reg_activation(reg_activation_14_4), .reg_weight(reg_weight_14_4), .reg_partial_sum(reg_psum_14_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_5( .activation_in(reg_activation_14_4), .weight_in(reg_weight_13_5), .partial_sum_in(reg_psum_13_5), .reg_activation(reg_activation_14_5), .reg_weight(reg_weight_14_5), .reg_partial_sum(reg_psum_14_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_6( .activation_in(reg_activation_14_5), .weight_in(reg_weight_13_6), .partial_sum_in(reg_psum_13_6), .reg_activation(reg_activation_14_6), .reg_weight(reg_weight_14_6), .reg_partial_sum(reg_psum_14_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_7( .activation_in(reg_activation_14_6), .weight_in(reg_weight_13_7), .partial_sum_in(reg_psum_13_7), .reg_activation(reg_activation_14_7), .reg_weight(reg_weight_14_7), .reg_partial_sum(reg_psum_14_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_8( .activation_in(reg_activation_14_7), .weight_in(reg_weight_13_8), .partial_sum_in(reg_psum_13_8), .reg_activation(reg_activation_14_8), .reg_weight(reg_weight_14_8), .reg_partial_sum(reg_psum_14_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_9( .activation_in(reg_activation_14_8), .weight_in(reg_weight_13_9), .partial_sum_in(reg_psum_13_9), .reg_activation(reg_activation_14_9), .reg_weight(reg_weight_14_9), .reg_partial_sum(reg_psum_14_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_10( .activation_in(reg_activation_14_9), .weight_in(reg_weight_13_10), .partial_sum_in(reg_psum_13_10), .reg_activation(reg_activation_14_10), .reg_weight(reg_weight_14_10), .reg_partial_sum(reg_psum_14_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_11( .activation_in(reg_activation_14_10), .weight_in(reg_weight_13_11), .partial_sum_in(reg_psum_13_11), .reg_activation(reg_activation_14_11), .reg_weight(reg_weight_14_11), .reg_partial_sum(reg_psum_14_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_12( .activation_in(reg_activation_14_11), .weight_in(reg_weight_13_12), .partial_sum_in(reg_psum_13_12), .reg_activation(reg_activation_14_12), .reg_weight(reg_weight_14_12), .reg_partial_sum(reg_psum_14_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_13( .activation_in(reg_activation_14_12), .weight_in(reg_weight_13_13), .partial_sum_in(reg_psum_13_13), .reg_activation(reg_activation_14_13), .reg_weight(reg_weight_14_13), .reg_partial_sum(reg_psum_14_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_14( .activation_in(reg_activation_14_13), .weight_in(reg_weight_13_14), .partial_sum_in(reg_psum_13_14), .reg_activation(reg_activation_14_14), .reg_weight(reg_weight_14_14), .reg_partial_sum(reg_psum_14_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_15( .activation_in(reg_activation_14_14), .weight_in(reg_weight_13_15), .partial_sum_in(reg_psum_13_15), .reg_activation(reg_activation_14_15), .reg_weight(reg_weight_14_15), .reg_partial_sum(reg_psum_14_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_16( .activation_in(reg_activation_14_15), .weight_in(reg_weight_13_16), .partial_sum_in(reg_psum_13_16), .reg_activation(reg_activation_14_16), .reg_weight(reg_weight_14_16), .reg_partial_sum(reg_psum_14_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_17( .activation_in(reg_activation_14_16), .weight_in(reg_weight_13_17), .partial_sum_in(reg_psum_13_17), .reg_activation(reg_activation_14_17), .reg_weight(reg_weight_14_17), .reg_partial_sum(reg_psum_14_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_18( .activation_in(reg_activation_14_17), .weight_in(reg_weight_13_18), .partial_sum_in(reg_psum_13_18), .reg_activation(reg_activation_14_18), .reg_weight(reg_weight_14_18), .reg_partial_sum(reg_psum_14_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_19( .activation_in(reg_activation_14_18), .weight_in(reg_weight_13_19), .partial_sum_in(reg_psum_13_19), .reg_activation(reg_activation_14_19), .reg_weight(reg_weight_14_19), .reg_partial_sum(reg_psum_14_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_20( .activation_in(reg_activation_14_19), .weight_in(reg_weight_13_20), .partial_sum_in(reg_psum_13_20), .reg_activation(reg_activation_14_20), .reg_weight(reg_weight_14_20), .reg_partial_sum(reg_psum_14_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_21( .activation_in(reg_activation_14_20), .weight_in(reg_weight_13_21), .partial_sum_in(reg_psum_13_21), .reg_activation(reg_activation_14_21), .reg_weight(reg_weight_14_21), .reg_partial_sum(reg_psum_14_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_22( .activation_in(reg_activation_14_21), .weight_in(reg_weight_13_22), .partial_sum_in(reg_psum_13_22), .reg_activation(reg_activation_14_22), .reg_weight(reg_weight_14_22), .reg_partial_sum(reg_psum_14_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_23( .activation_in(reg_activation_14_22), .weight_in(reg_weight_13_23), .partial_sum_in(reg_psum_13_23), .reg_activation(reg_activation_14_23), .reg_weight(reg_weight_14_23), .reg_partial_sum(reg_psum_14_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_24( .activation_in(reg_activation_14_23), .weight_in(reg_weight_13_24), .partial_sum_in(reg_psum_13_24), .reg_activation(reg_activation_14_24), .reg_weight(reg_weight_14_24), .reg_partial_sum(reg_psum_14_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_25( .activation_in(reg_activation_14_24), .weight_in(reg_weight_13_25), .partial_sum_in(reg_psum_13_25), .reg_activation(reg_activation_14_25), .reg_weight(reg_weight_14_25), .reg_partial_sum(reg_psum_14_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_26( .activation_in(reg_activation_14_25), .weight_in(reg_weight_13_26), .partial_sum_in(reg_psum_13_26), .reg_activation(reg_activation_14_26), .reg_weight(reg_weight_14_26), .reg_partial_sum(reg_psum_14_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_27( .activation_in(reg_activation_14_26), .weight_in(reg_weight_13_27), .partial_sum_in(reg_psum_13_27), .reg_activation(reg_activation_14_27), .reg_weight(reg_weight_14_27), .reg_partial_sum(reg_psum_14_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_28( .activation_in(reg_activation_14_27), .weight_in(reg_weight_13_28), .partial_sum_in(reg_psum_13_28), .reg_activation(reg_activation_14_28), .reg_weight(reg_weight_14_28), .reg_partial_sum(reg_psum_14_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_29( .activation_in(reg_activation_14_28), .weight_in(reg_weight_13_29), .partial_sum_in(reg_psum_13_29), .reg_activation(reg_activation_14_29), .reg_weight(reg_weight_14_29), .reg_partial_sum(reg_psum_14_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_30( .activation_in(reg_activation_14_29), .weight_in(reg_weight_13_30), .partial_sum_in(reg_psum_13_30), .reg_activation(reg_activation_14_30), .reg_weight(reg_weight_14_30), .reg_partial_sum(reg_psum_14_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_31( .activation_in(reg_activation_14_30), .weight_in(reg_weight_13_31), .partial_sum_in(reg_psum_13_31), .reg_activation(reg_activation_14_31), .reg_weight(reg_weight_14_31), .reg_partial_sum(reg_psum_14_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_32( .activation_in(reg_activation_14_31), .weight_in(reg_weight_13_32), .partial_sum_in(reg_psum_13_32), .reg_activation(reg_activation_14_32), .reg_weight(reg_weight_14_32), .reg_partial_sum(reg_psum_14_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_33( .activation_in(reg_activation_14_32), .weight_in(reg_weight_13_33), .partial_sum_in(reg_psum_13_33), .reg_activation(reg_activation_14_33), .reg_weight(reg_weight_14_33), .reg_partial_sum(reg_psum_14_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_34( .activation_in(reg_activation_14_33), .weight_in(reg_weight_13_34), .partial_sum_in(reg_psum_13_34), .reg_activation(reg_activation_14_34), .reg_weight(reg_weight_14_34), .reg_partial_sum(reg_psum_14_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_35( .activation_in(reg_activation_14_34), .weight_in(reg_weight_13_35), .partial_sum_in(reg_psum_13_35), .reg_activation(reg_activation_14_35), .reg_weight(reg_weight_14_35), .reg_partial_sum(reg_psum_14_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_36( .activation_in(reg_activation_14_35), .weight_in(reg_weight_13_36), .partial_sum_in(reg_psum_13_36), .reg_activation(reg_activation_14_36), .reg_weight(reg_weight_14_36), .reg_partial_sum(reg_psum_14_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_37( .activation_in(reg_activation_14_36), .weight_in(reg_weight_13_37), .partial_sum_in(reg_psum_13_37), .reg_activation(reg_activation_14_37), .reg_weight(reg_weight_14_37), .reg_partial_sum(reg_psum_14_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_38( .activation_in(reg_activation_14_37), .weight_in(reg_weight_13_38), .partial_sum_in(reg_psum_13_38), .reg_activation(reg_activation_14_38), .reg_weight(reg_weight_14_38), .reg_partial_sum(reg_psum_14_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_39( .activation_in(reg_activation_14_38), .weight_in(reg_weight_13_39), .partial_sum_in(reg_psum_13_39), .reg_activation(reg_activation_14_39), .reg_weight(reg_weight_14_39), .reg_partial_sum(reg_psum_14_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_40( .activation_in(reg_activation_14_39), .weight_in(reg_weight_13_40), .partial_sum_in(reg_psum_13_40), .reg_activation(reg_activation_14_40), .reg_weight(reg_weight_14_40), .reg_partial_sum(reg_psum_14_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_41( .activation_in(reg_activation_14_40), .weight_in(reg_weight_13_41), .partial_sum_in(reg_psum_13_41), .reg_activation(reg_activation_14_41), .reg_weight(reg_weight_14_41), .reg_partial_sum(reg_psum_14_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_42( .activation_in(reg_activation_14_41), .weight_in(reg_weight_13_42), .partial_sum_in(reg_psum_13_42), .reg_activation(reg_activation_14_42), .reg_weight(reg_weight_14_42), .reg_partial_sum(reg_psum_14_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_43( .activation_in(reg_activation_14_42), .weight_in(reg_weight_13_43), .partial_sum_in(reg_psum_13_43), .reg_activation(reg_activation_14_43), .reg_weight(reg_weight_14_43), .reg_partial_sum(reg_psum_14_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_44( .activation_in(reg_activation_14_43), .weight_in(reg_weight_13_44), .partial_sum_in(reg_psum_13_44), .reg_activation(reg_activation_14_44), .reg_weight(reg_weight_14_44), .reg_partial_sum(reg_psum_14_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_45( .activation_in(reg_activation_14_44), .weight_in(reg_weight_13_45), .partial_sum_in(reg_psum_13_45), .reg_activation(reg_activation_14_45), .reg_weight(reg_weight_14_45), .reg_partial_sum(reg_psum_14_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_46( .activation_in(reg_activation_14_45), .weight_in(reg_weight_13_46), .partial_sum_in(reg_psum_13_46), .reg_activation(reg_activation_14_46), .reg_weight(reg_weight_14_46), .reg_partial_sum(reg_psum_14_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_47( .activation_in(reg_activation_14_46), .weight_in(reg_weight_13_47), .partial_sum_in(reg_psum_13_47), .reg_activation(reg_activation_14_47), .reg_weight(reg_weight_14_47), .reg_partial_sum(reg_psum_14_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_48( .activation_in(reg_activation_14_47), .weight_in(reg_weight_13_48), .partial_sum_in(reg_psum_13_48), .reg_activation(reg_activation_14_48), .reg_weight(reg_weight_14_48), .reg_partial_sum(reg_psum_14_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_49( .activation_in(reg_activation_14_48), .weight_in(reg_weight_13_49), .partial_sum_in(reg_psum_13_49), .reg_activation(reg_activation_14_49), .reg_weight(reg_weight_14_49), .reg_partial_sum(reg_psum_14_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_50( .activation_in(reg_activation_14_49), .weight_in(reg_weight_13_50), .partial_sum_in(reg_psum_13_50), .reg_activation(reg_activation_14_50), .reg_weight(reg_weight_14_50), .reg_partial_sum(reg_psum_14_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_51( .activation_in(reg_activation_14_50), .weight_in(reg_weight_13_51), .partial_sum_in(reg_psum_13_51), .reg_activation(reg_activation_14_51), .reg_weight(reg_weight_14_51), .reg_partial_sum(reg_psum_14_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_52( .activation_in(reg_activation_14_51), .weight_in(reg_weight_13_52), .partial_sum_in(reg_psum_13_52), .reg_activation(reg_activation_14_52), .reg_weight(reg_weight_14_52), .reg_partial_sum(reg_psum_14_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_53( .activation_in(reg_activation_14_52), .weight_in(reg_weight_13_53), .partial_sum_in(reg_psum_13_53), .reg_activation(reg_activation_14_53), .reg_weight(reg_weight_14_53), .reg_partial_sum(reg_psum_14_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_54( .activation_in(reg_activation_14_53), .weight_in(reg_weight_13_54), .partial_sum_in(reg_psum_13_54), .reg_activation(reg_activation_14_54), .reg_weight(reg_weight_14_54), .reg_partial_sum(reg_psum_14_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_55( .activation_in(reg_activation_14_54), .weight_in(reg_weight_13_55), .partial_sum_in(reg_psum_13_55), .reg_activation(reg_activation_14_55), .reg_weight(reg_weight_14_55), .reg_partial_sum(reg_psum_14_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_56( .activation_in(reg_activation_14_55), .weight_in(reg_weight_13_56), .partial_sum_in(reg_psum_13_56), .reg_activation(reg_activation_14_56), .reg_weight(reg_weight_14_56), .reg_partial_sum(reg_psum_14_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_57( .activation_in(reg_activation_14_56), .weight_in(reg_weight_13_57), .partial_sum_in(reg_psum_13_57), .reg_activation(reg_activation_14_57), .reg_weight(reg_weight_14_57), .reg_partial_sum(reg_psum_14_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_58( .activation_in(reg_activation_14_57), .weight_in(reg_weight_13_58), .partial_sum_in(reg_psum_13_58), .reg_activation(reg_activation_14_58), .reg_weight(reg_weight_14_58), .reg_partial_sum(reg_psum_14_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_59( .activation_in(reg_activation_14_58), .weight_in(reg_weight_13_59), .partial_sum_in(reg_psum_13_59), .reg_activation(reg_activation_14_59), .reg_weight(reg_weight_14_59), .reg_partial_sum(reg_psum_14_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_60( .activation_in(reg_activation_14_59), .weight_in(reg_weight_13_60), .partial_sum_in(reg_psum_13_60), .reg_activation(reg_activation_14_60), .reg_weight(reg_weight_14_60), .reg_partial_sum(reg_psum_14_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_61( .activation_in(reg_activation_14_60), .weight_in(reg_weight_13_61), .partial_sum_in(reg_psum_13_61), .reg_activation(reg_activation_14_61), .reg_weight(reg_weight_14_61), .reg_partial_sum(reg_psum_14_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_62( .activation_in(reg_activation_14_61), .weight_in(reg_weight_13_62), .partial_sum_in(reg_psum_13_62), .reg_activation(reg_activation_14_62), .reg_weight(reg_weight_14_62), .reg_partial_sum(reg_psum_14_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_63( .activation_in(reg_activation_14_62), .weight_in(reg_weight_13_63), .partial_sum_in(reg_psum_13_63), .reg_weight(reg_weight_14_63), .reg_partial_sum(reg_psum_14_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_0( .activation_in(in_activation_15), .weight_in(reg_weight_14_0), .partial_sum_in(reg_psum_14_0), .reg_activation(reg_activation_15_0), .reg_weight(reg_weight_15_0), .reg_partial_sum(reg_psum_15_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_1( .activation_in(reg_activation_15_0), .weight_in(reg_weight_14_1), .partial_sum_in(reg_psum_14_1), .reg_activation(reg_activation_15_1), .reg_weight(reg_weight_15_1), .reg_partial_sum(reg_psum_15_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_2( .activation_in(reg_activation_15_1), .weight_in(reg_weight_14_2), .partial_sum_in(reg_psum_14_2), .reg_activation(reg_activation_15_2), .reg_weight(reg_weight_15_2), .reg_partial_sum(reg_psum_15_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_3( .activation_in(reg_activation_15_2), .weight_in(reg_weight_14_3), .partial_sum_in(reg_psum_14_3), .reg_activation(reg_activation_15_3), .reg_weight(reg_weight_15_3), .reg_partial_sum(reg_psum_15_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_4( .activation_in(reg_activation_15_3), .weight_in(reg_weight_14_4), .partial_sum_in(reg_psum_14_4), .reg_activation(reg_activation_15_4), .reg_weight(reg_weight_15_4), .reg_partial_sum(reg_psum_15_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_5( .activation_in(reg_activation_15_4), .weight_in(reg_weight_14_5), .partial_sum_in(reg_psum_14_5), .reg_activation(reg_activation_15_5), .reg_weight(reg_weight_15_5), .reg_partial_sum(reg_psum_15_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_6( .activation_in(reg_activation_15_5), .weight_in(reg_weight_14_6), .partial_sum_in(reg_psum_14_6), .reg_activation(reg_activation_15_6), .reg_weight(reg_weight_15_6), .reg_partial_sum(reg_psum_15_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_7( .activation_in(reg_activation_15_6), .weight_in(reg_weight_14_7), .partial_sum_in(reg_psum_14_7), .reg_activation(reg_activation_15_7), .reg_weight(reg_weight_15_7), .reg_partial_sum(reg_psum_15_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_8( .activation_in(reg_activation_15_7), .weight_in(reg_weight_14_8), .partial_sum_in(reg_psum_14_8), .reg_activation(reg_activation_15_8), .reg_weight(reg_weight_15_8), .reg_partial_sum(reg_psum_15_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_9( .activation_in(reg_activation_15_8), .weight_in(reg_weight_14_9), .partial_sum_in(reg_psum_14_9), .reg_activation(reg_activation_15_9), .reg_weight(reg_weight_15_9), .reg_partial_sum(reg_psum_15_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_10( .activation_in(reg_activation_15_9), .weight_in(reg_weight_14_10), .partial_sum_in(reg_psum_14_10), .reg_activation(reg_activation_15_10), .reg_weight(reg_weight_15_10), .reg_partial_sum(reg_psum_15_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_11( .activation_in(reg_activation_15_10), .weight_in(reg_weight_14_11), .partial_sum_in(reg_psum_14_11), .reg_activation(reg_activation_15_11), .reg_weight(reg_weight_15_11), .reg_partial_sum(reg_psum_15_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_12( .activation_in(reg_activation_15_11), .weight_in(reg_weight_14_12), .partial_sum_in(reg_psum_14_12), .reg_activation(reg_activation_15_12), .reg_weight(reg_weight_15_12), .reg_partial_sum(reg_psum_15_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_13( .activation_in(reg_activation_15_12), .weight_in(reg_weight_14_13), .partial_sum_in(reg_psum_14_13), .reg_activation(reg_activation_15_13), .reg_weight(reg_weight_15_13), .reg_partial_sum(reg_psum_15_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_14( .activation_in(reg_activation_15_13), .weight_in(reg_weight_14_14), .partial_sum_in(reg_psum_14_14), .reg_activation(reg_activation_15_14), .reg_weight(reg_weight_15_14), .reg_partial_sum(reg_psum_15_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_15( .activation_in(reg_activation_15_14), .weight_in(reg_weight_14_15), .partial_sum_in(reg_psum_14_15), .reg_activation(reg_activation_15_15), .reg_weight(reg_weight_15_15), .reg_partial_sum(reg_psum_15_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_16( .activation_in(reg_activation_15_15), .weight_in(reg_weight_14_16), .partial_sum_in(reg_psum_14_16), .reg_activation(reg_activation_15_16), .reg_weight(reg_weight_15_16), .reg_partial_sum(reg_psum_15_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_17( .activation_in(reg_activation_15_16), .weight_in(reg_weight_14_17), .partial_sum_in(reg_psum_14_17), .reg_activation(reg_activation_15_17), .reg_weight(reg_weight_15_17), .reg_partial_sum(reg_psum_15_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_18( .activation_in(reg_activation_15_17), .weight_in(reg_weight_14_18), .partial_sum_in(reg_psum_14_18), .reg_activation(reg_activation_15_18), .reg_weight(reg_weight_15_18), .reg_partial_sum(reg_psum_15_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_19( .activation_in(reg_activation_15_18), .weight_in(reg_weight_14_19), .partial_sum_in(reg_psum_14_19), .reg_activation(reg_activation_15_19), .reg_weight(reg_weight_15_19), .reg_partial_sum(reg_psum_15_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_20( .activation_in(reg_activation_15_19), .weight_in(reg_weight_14_20), .partial_sum_in(reg_psum_14_20), .reg_activation(reg_activation_15_20), .reg_weight(reg_weight_15_20), .reg_partial_sum(reg_psum_15_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_21( .activation_in(reg_activation_15_20), .weight_in(reg_weight_14_21), .partial_sum_in(reg_psum_14_21), .reg_activation(reg_activation_15_21), .reg_weight(reg_weight_15_21), .reg_partial_sum(reg_psum_15_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_22( .activation_in(reg_activation_15_21), .weight_in(reg_weight_14_22), .partial_sum_in(reg_psum_14_22), .reg_activation(reg_activation_15_22), .reg_weight(reg_weight_15_22), .reg_partial_sum(reg_psum_15_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_23( .activation_in(reg_activation_15_22), .weight_in(reg_weight_14_23), .partial_sum_in(reg_psum_14_23), .reg_activation(reg_activation_15_23), .reg_weight(reg_weight_15_23), .reg_partial_sum(reg_psum_15_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_24( .activation_in(reg_activation_15_23), .weight_in(reg_weight_14_24), .partial_sum_in(reg_psum_14_24), .reg_activation(reg_activation_15_24), .reg_weight(reg_weight_15_24), .reg_partial_sum(reg_psum_15_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_25( .activation_in(reg_activation_15_24), .weight_in(reg_weight_14_25), .partial_sum_in(reg_psum_14_25), .reg_activation(reg_activation_15_25), .reg_weight(reg_weight_15_25), .reg_partial_sum(reg_psum_15_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_26( .activation_in(reg_activation_15_25), .weight_in(reg_weight_14_26), .partial_sum_in(reg_psum_14_26), .reg_activation(reg_activation_15_26), .reg_weight(reg_weight_15_26), .reg_partial_sum(reg_psum_15_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_27( .activation_in(reg_activation_15_26), .weight_in(reg_weight_14_27), .partial_sum_in(reg_psum_14_27), .reg_activation(reg_activation_15_27), .reg_weight(reg_weight_15_27), .reg_partial_sum(reg_psum_15_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_28( .activation_in(reg_activation_15_27), .weight_in(reg_weight_14_28), .partial_sum_in(reg_psum_14_28), .reg_activation(reg_activation_15_28), .reg_weight(reg_weight_15_28), .reg_partial_sum(reg_psum_15_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_29( .activation_in(reg_activation_15_28), .weight_in(reg_weight_14_29), .partial_sum_in(reg_psum_14_29), .reg_activation(reg_activation_15_29), .reg_weight(reg_weight_15_29), .reg_partial_sum(reg_psum_15_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_30( .activation_in(reg_activation_15_29), .weight_in(reg_weight_14_30), .partial_sum_in(reg_psum_14_30), .reg_activation(reg_activation_15_30), .reg_weight(reg_weight_15_30), .reg_partial_sum(reg_psum_15_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_31( .activation_in(reg_activation_15_30), .weight_in(reg_weight_14_31), .partial_sum_in(reg_psum_14_31), .reg_activation(reg_activation_15_31), .reg_weight(reg_weight_15_31), .reg_partial_sum(reg_psum_15_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_32( .activation_in(reg_activation_15_31), .weight_in(reg_weight_14_32), .partial_sum_in(reg_psum_14_32), .reg_activation(reg_activation_15_32), .reg_weight(reg_weight_15_32), .reg_partial_sum(reg_psum_15_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_33( .activation_in(reg_activation_15_32), .weight_in(reg_weight_14_33), .partial_sum_in(reg_psum_14_33), .reg_activation(reg_activation_15_33), .reg_weight(reg_weight_15_33), .reg_partial_sum(reg_psum_15_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_34( .activation_in(reg_activation_15_33), .weight_in(reg_weight_14_34), .partial_sum_in(reg_psum_14_34), .reg_activation(reg_activation_15_34), .reg_weight(reg_weight_15_34), .reg_partial_sum(reg_psum_15_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_35( .activation_in(reg_activation_15_34), .weight_in(reg_weight_14_35), .partial_sum_in(reg_psum_14_35), .reg_activation(reg_activation_15_35), .reg_weight(reg_weight_15_35), .reg_partial_sum(reg_psum_15_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_36( .activation_in(reg_activation_15_35), .weight_in(reg_weight_14_36), .partial_sum_in(reg_psum_14_36), .reg_activation(reg_activation_15_36), .reg_weight(reg_weight_15_36), .reg_partial_sum(reg_psum_15_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_37( .activation_in(reg_activation_15_36), .weight_in(reg_weight_14_37), .partial_sum_in(reg_psum_14_37), .reg_activation(reg_activation_15_37), .reg_weight(reg_weight_15_37), .reg_partial_sum(reg_psum_15_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_38( .activation_in(reg_activation_15_37), .weight_in(reg_weight_14_38), .partial_sum_in(reg_psum_14_38), .reg_activation(reg_activation_15_38), .reg_weight(reg_weight_15_38), .reg_partial_sum(reg_psum_15_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_39( .activation_in(reg_activation_15_38), .weight_in(reg_weight_14_39), .partial_sum_in(reg_psum_14_39), .reg_activation(reg_activation_15_39), .reg_weight(reg_weight_15_39), .reg_partial_sum(reg_psum_15_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_40( .activation_in(reg_activation_15_39), .weight_in(reg_weight_14_40), .partial_sum_in(reg_psum_14_40), .reg_activation(reg_activation_15_40), .reg_weight(reg_weight_15_40), .reg_partial_sum(reg_psum_15_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_41( .activation_in(reg_activation_15_40), .weight_in(reg_weight_14_41), .partial_sum_in(reg_psum_14_41), .reg_activation(reg_activation_15_41), .reg_weight(reg_weight_15_41), .reg_partial_sum(reg_psum_15_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_42( .activation_in(reg_activation_15_41), .weight_in(reg_weight_14_42), .partial_sum_in(reg_psum_14_42), .reg_activation(reg_activation_15_42), .reg_weight(reg_weight_15_42), .reg_partial_sum(reg_psum_15_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_43( .activation_in(reg_activation_15_42), .weight_in(reg_weight_14_43), .partial_sum_in(reg_psum_14_43), .reg_activation(reg_activation_15_43), .reg_weight(reg_weight_15_43), .reg_partial_sum(reg_psum_15_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_44( .activation_in(reg_activation_15_43), .weight_in(reg_weight_14_44), .partial_sum_in(reg_psum_14_44), .reg_activation(reg_activation_15_44), .reg_weight(reg_weight_15_44), .reg_partial_sum(reg_psum_15_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_45( .activation_in(reg_activation_15_44), .weight_in(reg_weight_14_45), .partial_sum_in(reg_psum_14_45), .reg_activation(reg_activation_15_45), .reg_weight(reg_weight_15_45), .reg_partial_sum(reg_psum_15_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_46( .activation_in(reg_activation_15_45), .weight_in(reg_weight_14_46), .partial_sum_in(reg_psum_14_46), .reg_activation(reg_activation_15_46), .reg_weight(reg_weight_15_46), .reg_partial_sum(reg_psum_15_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_47( .activation_in(reg_activation_15_46), .weight_in(reg_weight_14_47), .partial_sum_in(reg_psum_14_47), .reg_activation(reg_activation_15_47), .reg_weight(reg_weight_15_47), .reg_partial_sum(reg_psum_15_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_48( .activation_in(reg_activation_15_47), .weight_in(reg_weight_14_48), .partial_sum_in(reg_psum_14_48), .reg_activation(reg_activation_15_48), .reg_weight(reg_weight_15_48), .reg_partial_sum(reg_psum_15_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_49( .activation_in(reg_activation_15_48), .weight_in(reg_weight_14_49), .partial_sum_in(reg_psum_14_49), .reg_activation(reg_activation_15_49), .reg_weight(reg_weight_15_49), .reg_partial_sum(reg_psum_15_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_50( .activation_in(reg_activation_15_49), .weight_in(reg_weight_14_50), .partial_sum_in(reg_psum_14_50), .reg_activation(reg_activation_15_50), .reg_weight(reg_weight_15_50), .reg_partial_sum(reg_psum_15_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_51( .activation_in(reg_activation_15_50), .weight_in(reg_weight_14_51), .partial_sum_in(reg_psum_14_51), .reg_activation(reg_activation_15_51), .reg_weight(reg_weight_15_51), .reg_partial_sum(reg_psum_15_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_52( .activation_in(reg_activation_15_51), .weight_in(reg_weight_14_52), .partial_sum_in(reg_psum_14_52), .reg_activation(reg_activation_15_52), .reg_weight(reg_weight_15_52), .reg_partial_sum(reg_psum_15_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_53( .activation_in(reg_activation_15_52), .weight_in(reg_weight_14_53), .partial_sum_in(reg_psum_14_53), .reg_activation(reg_activation_15_53), .reg_weight(reg_weight_15_53), .reg_partial_sum(reg_psum_15_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_54( .activation_in(reg_activation_15_53), .weight_in(reg_weight_14_54), .partial_sum_in(reg_psum_14_54), .reg_activation(reg_activation_15_54), .reg_weight(reg_weight_15_54), .reg_partial_sum(reg_psum_15_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_55( .activation_in(reg_activation_15_54), .weight_in(reg_weight_14_55), .partial_sum_in(reg_psum_14_55), .reg_activation(reg_activation_15_55), .reg_weight(reg_weight_15_55), .reg_partial_sum(reg_psum_15_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_56( .activation_in(reg_activation_15_55), .weight_in(reg_weight_14_56), .partial_sum_in(reg_psum_14_56), .reg_activation(reg_activation_15_56), .reg_weight(reg_weight_15_56), .reg_partial_sum(reg_psum_15_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_57( .activation_in(reg_activation_15_56), .weight_in(reg_weight_14_57), .partial_sum_in(reg_psum_14_57), .reg_activation(reg_activation_15_57), .reg_weight(reg_weight_15_57), .reg_partial_sum(reg_psum_15_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_58( .activation_in(reg_activation_15_57), .weight_in(reg_weight_14_58), .partial_sum_in(reg_psum_14_58), .reg_activation(reg_activation_15_58), .reg_weight(reg_weight_15_58), .reg_partial_sum(reg_psum_15_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_59( .activation_in(reg_activation_15_58), .weight_in(reg_weight_14_59), .partial_sum_in(reg_psum_14_59), .reg_activation(reg_activation_15_59), .reg_weight(reg_weight_15_59), .reg_partial_sum(reg_psum_15_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_60( .activation_in(reg_activation_15_59), .weight_in(reg_weight_14_60), .partial_sum_in(reg_psum_14_60), .reg_activation(reg_activation_15_60), .reg_weight(reg_weight_15_60), .reg_partial_sum(reg_psum_15_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_61( .activation_in(reg_activation_15_60), .weight_in(reg_weight_14_61), .partial_sum_in(reg_psum_14_61), .reg_activation(reg_activation_15_61), .reg_weight(reg_weight_15_61), .reg_partial_sum(reg_psum_15_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_62( .activation_in(reg_activation_15_61), .weight_in(reg_weight_14_62), .partial_sum_in(reg_psum_14_62), .reg_activation(reg_activation_15_62), .reg_weight(reg_weight_15_62), .reg_partial_sum(reg_psum_15_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_63( .activation_in(reg_activation_15_62), .weight_in(reg_weight_14_63), .partial_sum_in(reg_psum_14_63), .reg_weight(reg_weight_15_63), .reg_partial_sum(reg_psum_15_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_0( .activation_in(in_activation_16), .weight_in(reg_weight_15_0), .partial_sum_in(reg_psum_15_0), .reg_activation(reg_activation_16_0), .reg_weight(reg_weight_16_0), .reg_partial_sum(reg_psum_16_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_1( .activation_in(reg_activation_16_0), .weight_in(reg_weight_15_1), .partial_sum_in(reg_psum_15_1), .reg_activation(reg_activation_16_1), .reg_weight(reg_weight_16_1), .reg_partial_sum(reg_psum_16_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_2( .activation_in(reg_activation_16_1), .weight_in(reg_weight_15_2), .partial_sum_in(reg_psum_15_2), .reg_activation(reg_activation_16_2), .reg_weight(reg_weight_16_2), .reg_partial_sum(reg_psum_16_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_3( .activation_in(reg_activation_16_2), .weight_in(reg_weight_15_3), .partial_sum_in(reg_psum_15_3), .reg_activation(reg_activation_16_3), .reg_weight(reg_weight_16_3), .reg_partial_sum(reg_psum_16_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_4( .activation_in(reg_activation_16_3), .weight_in(reg_weight_15_4), .partial_sum_in(reg_psum_15_4), .reg_activation(reg_activation_16_4), .reg_weight(reg_weight_16_4), .reg_partial_sum(reg_psum_16_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_5( .activation_in(reg_activation_16_4), .weight_in(reg_weight_15_5), .partial_sum_in(reg_psum_15_5), .reg_activation(reg_activation_16_5), .reg_weight(reg_weight_16_5), .reg_partial_sum(reg_psum_16_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_6( .activation_in(reg_activation_16_5), .weight_in(reg_weight_15_6), .partial_sum_in(reg_psum_15_6), .reg_activation(reg_activation_16_6), .reg_weight(reg_weight_16_6), .reg_partial_sum(reg_psum_16_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_7( .activation_in(reg_activation_16_6), .weight_in(reg_weight_15_7), .partial_sum_in(reg_psum_15_7), .reg_activation(reg_activation_16_7), .reg_weight(reg_weight_16_7), .reg_partial_sum(reg_psum_16_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_8( .activation_in(reg_activation_16_7), .weight_in(reg_weight_15_8), .partial_sum_in(reg_psum_15_8), .reg_activation(reg_activation_16_8), .reg_weight(reg_weight_16_8), .reg_partial_sum(reg_psum_16_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_9( .activation_in(reg_activation_16_8), .weight_in(reg_weight_15_9), .partial_sum_in(reg_psum_15_9), .reg_activation(reg_activation_16_9), .reg_weight(reg_weight_16_9), .reg_partial_sum(reg_psum_16_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_10( .activation_in(reg_activation_16_9), .weight_in(reg_weight_15_10), .partial_sum_in(reg_psum_15_10), .reg_activation(reg_activation_16_10), .reg_weight(reg_weight_16_10), .reg_partial_sum(reg_psum_16_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_11( .activation_in(reg_activation_16_10), .weight_in(reg_weight_15_11), .partial_sum_in(reg_psum_15_11), .reg_activation(reg_activation_16_11), .reg_weight(reg_weight_16_11), .reg_partial_sum(reg_psum_16_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_12( .activation_in(reg_activation_16_11), .weight_in(reg_weight_15_12), .partial_sum_in(reg_psum_15_12), .reg_activation(reg_activation_16_12), .reg_weight(reg_weight_16_12), .reg_partial_sum(reg_psum_16_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_13( .activation_in(reg_activation_16_12), .weight_in(reg_weight_15_13), .partial_sum_in(reg_psum_15_13), .reg_activation(reg_activation_16_13), .reg_weight(reg_weight_16_13), .reg_partial_sum(reg_psum_16_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_14( .activation_in(reg_activation_16_13), .weight_in(reg_weight_15_14), .partial_sum_in(reg_psum_15_14), .reg_activation(reg_activation_16_14), .reg_weight(reg_weight_16_14), .reg_partial_sum(reg_psum_16_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_15( .activation_in(reg_activation_16_14), .weight_in(reg_weight_15_15), .partial_sum_in(reg_psum_15_15), .reg_activation(reg_activation_16_15), .reg_weight(reg_weight_16_15), .reg_partial_sum(reg_psum_16_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_16( .activation_in(reg_activation_16_15), .weight_in(reg_weight_15_16), .partial_sum_in(reg_psum_15_16), .reg_activation(reg_activation_16_16), .reg_weight(reg_weight_16_16), .reg_partial_sum(reg_psum_16_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_17( .activation_in(reg_activation_16_16), .weight_in(reg_weight_15_17), .partial_sum_in(reg_psum_15_17), .reg_activation(reg_activation_16_17), .reg_weight(reg_weight_16_17), .reg_partial_sum(reg_psum_16_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_18( .activation_in(reg_activation_16_17), .weight_in(reg_weight_15_18), .partial_sum_in(reg_psum_15_18), .reg_activation(reg_activation_16_18), .reg_weight(reg_weight_16_18), .reg_partial_sum(reg_psum_16_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_19( .activation_in(reg_activation_16_18), .weight_in(reg_weight_15_19), .partial_sum_in(reg_psum_15_19), .reg_activation(reg_activation_16_19), .reg_weight(reg_weight_16_19), .reg_partial_sum(reg_psum_16_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_20( .activation_in(reg_activation_16_19), .weight_in(reg_weight_15_20), .partial_sum_in(reg_psum_15_20), .reg_activation(reg_activation_16_20), .reg_weight(reg_weight_16_20), .reg_partial_sum(reg_psum_16_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_21( .activation_in(reg_activation_16_20), .weight_in(reg_weight_15_21), .partial_sum_in(reg_psum_15_21), .reg_activation(reg_activation_16_21), .reg_weight(reg_weight_16_21), .reg_partial_sum(reg_psum_16_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_22( .activation_in(reg_activation_16_21), .weight_in(reg_weight_15_22), .partial_sum_in(reg_psum_15_22), .reg_activation(reg_activation_16_22), .reg_weight(reg_weight_16_22), .reg_partial_sum(reg_psum_16_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_23( .activation_in(reg_activation_16_22), .weight_in(reg_weight_15_23), .partial_sum_in(reg_psum_15_23), .reg_activation(reg_activation_16_23), .reg_weight(reg_weight_16_23), .reg_partial_sum(reg_psum_16_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_24( .activation_in(reg_activation_16_23), .weight_in(reg_weight_15_24), .partial_sum_in(reg_psum_15_24), .reg_activation(reg_activation_16_24), .reg_weight(reg_weight_16_24), .reg_partial_sum(reg_psum_16_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_25( .activation_in(reg_activation_16_24), .weight_in(reg_weight_15_25), .partial_sum_in(reg_psum_15_25), .reg_activation(reg_activation_16_25), .reg_weight(reg_weight_16_25), .reg_partial_sum(reg_psum_16_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_26( .activation_in(reg_activation_16_25), .weight_in(reg_weight_15_26), .partial_sum_in(reg_psum_15_26), .reg_activation(reg_activation_16_26), .reg_weight(reg_weight_16_26), .reg_partial_sum(reg_psum_16_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_27( .activation_in(reg_activation_16_26), .weight_in(reg_weight_15_27), .partial_sum_in(reg_psum_15_27), .reg_activation(reg_activation_16_27), .reg_weight(reg_weight_16_27), .reg_partial_sum(reg_psum_16_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_28( .activation_in(reg_activation_16_27), .weight_in(reg_weight_15_28), .partial_sum_in(reg_psum_15_28), .reg_activation(reg_activation_16_28), .reg_weight(reg_weight_16_28), .reg_partial_sum(reg_psum_16_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_29( .activation_in(reg_activation_16_28), .weight_in(reg_weight_15_29), .partial_sum_in(reg_psum_15_29), .reg_activation(reg_activation_16_29), .reg_weight(reg_weight_16_29), .reg_partial_sum(reg_psum_16_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_30( .activation_in(reg_activation_16_29), .weight_in(reg_weight_15_30), .partial_sum_in(reg_psum_15_30), .reg_activation(reg_activation_16_30), .reg_weight(reg_weight_16_30), .reg_partial_sum(reg_psum_16_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_31( .activation_in(reg_activation_16_30), .weight_in(reg_weight_15_31), .partial_sum_in(reg_psum_15_31), .reg_activation(reg_activation_16_31), .reg_weight(reg_weight_16_31), .reg_partial_sum(reg_psum_16_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_32( .activation_in(reg_activation_16_31), .weight_in(reg_weight_15_32), .partial_sum_in(reg_psum_15_32), .reg_activation(reg_activation_16_32), .reg_weight(reg_weight_16_32), .reg_partial_sum(reg_psum_16_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_33( .activation_in(reg_activation_16_32), .weight_in(reg_weight_15_33), .partial_sum_in(reg_psum_15_33), .reg_activation(reg_activation_16_33), .reg_weight(reg_weight_16_33), .reg_partial_sum(reg_psum_16_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_34( .activation_in(reg_activation_16_33), .weight_in(reg_weight_15_34), .partial_sum_in(reg_psum_15_34), .reg_activation(reg_activation_16_34), .reg_weight(reg_weight_16_34), .reg_partial_sum(reg_psum_16_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_35( .activation_in(reg_activation_16_34), .weight_in(reg_weight_15_35), .partial_sum_in(reg_psum_15_35), .reg_activation(reg_activation_16_35), .reg_weight(reg_weight_16_35), .reg_partial_sum(reg_psum_16_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_36( .activation_in(reg_activation_16_35), .weight_in(reg_weight_15_36), .partial_sum_in(reg_psum_15_36), .reg_activation(reg_activation_16_36), .reg_weight(reg_weight_16_36), .reg_partial_sum(reg_psum_16_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_37( .activation_in(reg_activation_16_36), .weight_in(reg_weight_15_37), .partial_sum_in(reg_psum_15_37), .reg_activation(reg_activation_16_37), .reg_weight(reg_weight_16_37), .reg_partial_sum(reg_psum_16_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_38( .activation_in(reg_activation_16_37), .weight_in(reg_weight_15_38), .partial_sum_in(reg_psum_15_38), .reg_activation(reg_activation_16_38), .reg_weight(reg_weight_16_38), .reg_partial_sum(reg_psum_16_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_39( .activation_in(reg_activation_16_38), .weight_in(reg_weight_15_39), .partial_sum_in(reg_psum_15_39), .reg_activation(reg_activation_16_39), .reg_weight(reg_weight_16_39), .reg_partial_sum(reg_psum_16_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_40( .activation_in(reg_activation_16_39), .weight_in(reg_weight_15_40), .partial_sum_in(reg_psum_15_40), .reg_activation(reg_activation_16_40), .reg_weight(reg_weight_16_40), .reg_partial_sum(reg_psum_16_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_41( .activation_in(reg_activation_16_40), .weight_in(reg_weight_15_41), .partial_sum_in(reg_psum_15_41), .reg_activation(reg_activation_16_41), .reg_weight(reg_weight_16_41), .reg_partial_sum(reg_psum_16_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_42( .activation_in(reg_activation_16_41), .weight_in(reg_weight_15_42), .partial_sum_in(reg_psum_15_42), .reg_activation(reg_activation_16_42), .reg_weight(reg_weight_16_42), .reg_partial_sum(reg_psum_16_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_43( .activation_in(reg_activation_16_42), .weight_in(reg_weight_15_43), .partial_sum_in(reg_psum_15_43), .reg_activation(reg_activation_16_43), .reg_weight(reg_weight_16_43), .reg_partial_sum(reg_psum_16_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_44( .activation_in(reg_activation_16_43), .weight_in(reg_weight_15_44), .partial_sum_in(reg_psum_15_44), .reg_activation(reg_activation_16_44), .reg_weight(reg_weight_16_44), .reg_partial_sum(reg_psum_16_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_45( .activation_in(reg_activation_16_44), .weight_in(reg_weight_15_45), .partial_sum_in(reg_psum_15_45), .reg_activation(reg_activation_16_45), .reg_weight(reg_weight_16_45), .reg_partial_sum(reg_psum_16_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_46( .activation_in(reg_activation_16_45), .weight_in(reg_weight_15_46), .partial_sum_in(reg_psum_15_46), .reg_activation(reg_activation_16_46), .reg_weight(reg_weight_16_46), .reg_partial_sum(reg_psum_16_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_47( .activation_in(reg_activation_16_46), .weight_in(reg_weight_15_47), .partial_sum_in(reg_psum_15_47), .reg_activation(reg_activation_16_47), .reg_weight(reg_weight_16_47), .reg_partial_sum(reg_psum_16_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_48( .activation_in(reg_activation_16_47), .weight_in(reg_weight_15_48), .partial_sum_in(reg_psum_15_48), .reg_activation(reg_activation_16_48), .reg_weight(reg_weight_16_48), .reg_partial_sum(reg_psum_16_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_49( .activation_in(reg_activation_16_48), .weight_in(reg_weight_15_49), .partial_sum_in(reg_psum_15_49), .reg_activation(reg_activation_16_49), .reg_weight(reg_weight_16_49), .reg_partial_sum(reg_psum_16_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_50( .activation_in(reg_activation_16_49), .weight_in(reg_weight_15_50), .partial_sum_in(reg_psum_15_50), .reg_activation(reg_activation_16_50), .reg_weight(reg_weight_16_50), .reg_partial_sum(reg_psum_16_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_51( .activation_in(reg_activation_16_50), .weight_in(reg_weight_15_51), .partial_sum_in(reg_psum_15_51), .reg_activation(reg_activation_16_51), .reg_weight(reg_weight_16_51), .reg_partial_sum(reg_psum_16_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_52( .activation_in(reg_activation_16_51), .weight_in(reg_weight_15_52), .partial_sum_in(reg_psum_15_52), .reg_activation(reg_activation_16_52), .reg_weight(reg_weight_16_52), .reg_partial_sum(reg_psum_16_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_53( .activation_in(reg_activation_16_52), .weight_in(reg_weight_15_53), .partial_sum_in(reg_psum_15_53), .reg_activation(reg_activation_16_53), .reg_weight(reg_weight_16_53), .reg_partial_sum(reg_psum_16_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_54( .activation_in(reg_activation_16_53), .weight_in(reg_weight_15_54), .partial_sum_in(reg_psum_15_54), .reg_activation(reg_activation_16_54), .reg_weight(reg_weight_16_54), .reg_partial_sum(reg_psum_16_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_55( .activation_in(reg_activation_16_54), .weight_in(reg_weight_15_55), .partial_sum_in(reg_psum_15_55), .reg_activation(reg_activation_16_55), .reg_weight(reg_weight_16_55), .reg_partial_sum(reg_psum_16_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_56( .activation_in(reg_activation_16_55), .weight_in(reg_weight_15_56), .partial_sum_in(reg_psum_15_56), .reg_activation(reg_activation_16_56), .reg_weight(reg_weight_16_56), .reg_partial_sum(reg_psum_16_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_57( .activation_in(reg_activation_16_56), .weight_in(reg_weight_15_57), .partial_sum_in(reg_psum_15_57), .reg_activation(reg_activation_16_57), .reg_weight(reg_weight_16_57), .reg_partial_sum(reg_psum_16_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_58( .activation_in(reg_activation_16_57), .weight_in(reg_weight_15_58), .partial_sum_in(reg_psum_15_58), .reg_activation(reg_activation_16_58), .reg_weight(reg_weight_16_58), .reg_partial_sum(reg_psum_16_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_59( .activation_in(reg_activation_16_58), .weight_in(reg_weight_15_59), .partial_sum_in(reg_psum_15_59), .reg_activation(reg_activation_16_59), .reg_weight(reg_weight_16_59), .reg_partial_sum(reg_psum_16_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_60( .activation_in(reg_activation_16_59), .weight_in(reg_weight_15_60), .partial_sum_in(reg_psum_15_60), .reg_activation(reg_activation_16_60), .reg_weight(reg_weight_16_60), .reg_partial_sum(reg_psum_16_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_61( .activation_in(reg_activation_16_60), .weight_in(reg_weight_15_61), .partial_sum_in(reg_psum_15_61), .reg_activation(reg_activation_16_61), .reg_weight(reg_weight_16_61), .reg_partial_sum(reg_psum_16_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_62( .activation_in(reg_activation_16_61), .weight_in(reg_weight_15_62), .partial_sum_in(reg_psum_15_62), .reg_activation(reg_activation_16_62), .reg_weight(reg_weight_16_62), .reg_partial_sum(reg_psum_16_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_63( .activation_in(reg_activation_16_62), .weight_in(reg_weight_15_63), .partial_sum_in(reg_psum_15_63), .reg_weight(reg_weight_16_63), .reg_partial_sum(reg_psum_16_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_0( .activation_in(in_activation_17), .weight_in(reg_weight_16_0), .partial_sum_in(reg_psum_16_0), .reg_activation(reg_activation_17_0), .reg_weight(reg_weight_17_0), .reg_partial_sum(reg_psum_17_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_1( .activation_in(reg_activation_17_0), .weight_in(reg_weight_16_1), .partial_sum_in(reg_psum_16_1), .reg_activation(reg_activation_17_1), .reg_weight(reg_weight_17_1), .reg_partial_sum(reg_psum_17_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_2( .activation_in(reg_activation_17_1), .weight_in(reg_weight_16_2), .partial_sum_in(reg_psum_16_2), .reg_activation(reg_activation_17_2), .reg_weight(reg_weight_17_2), .reg_partial_sum(reg_psum_17_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_3( .activation_in(reg_activation_17_2), .weight_in(reg_weight_16_3), .partial_sum_in(reg_psum_16_3), .reg_activation(reg_activation_17_3), .reg_weight(reg_weight_17_3), .reg_partial_sum(reg_psum_17_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_4( .activation_in(reg_activation_17_3), .weight_in(reg_weight_16_4), .partial_sum_in(reg_psum_16_4), .reg_activation(reg_activation_17_4), .reg_weight(reg_weight_17_4), .reg_partial_sum(reg_psum_17_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_5( .activation_in(reg_activation_17_4), .weight_in(reg_weight_16_5), .partial_sum_in(reg_psum_16_5), .reg_activation(reg_activation_17_5), .reg_weight(reg_weight_17_5), .reg_partial_sum(reg_psum_17_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_6( .activation_in(reg_activation_17_5), .weight_in(reg_weight_16_6), .partial_sum_in(reg_psum_16_6), .reg_activation(reg_activation_17_6), .reg_weight(reg_weight_17_6), .reg_partial_sum(reg_psum_17_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_7( .activation_in(reg_activation_17_6), .weight_in(reg_weight_16_7), .partial_sum_in(reg_psum_16_7), .reg_activation(reg_activation_17_7), .reg_weight(reg_weight_17_7), .reg_partial_sum(reg_psum_17_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_8( .activation_in(reg_activation_17_7), .weight_in(reg_weight_16_8), .partial_sum_in(reg_psum_16_8), .reg_activation(reg_activation_17_8), .reg_weight(reg_weight_17_8), .reg_partial_sum(reg_psum_17_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_9( .activation_in(reg_activation_17_8), .weight_in(reg_weight_16_9), .partial_sum_in(reg_psum_16_9), .reg_activation(reg_activation_17_9), .reg_weight(reg_weight_17_9), .reg_partial_sum(reg_psum_17_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_10( .activation_in(reg_activation_17_9), .weight_in(reg_weight_16_10), .partial_sum_in(reg_psum_16_10), .reg_activation(reg_activation_17_10), .reg_weight(reg_weight_17_10), .reg_partial_sum(reg_psum_17_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_11( .activation_in(reg_activation_17_10), .weight_in(reg_weight_16_11), .partial_sum_in(reg_psum_16_11), .reg_activation(reg_activation_17_11), .reg_weight(reg_weight_17_11), .reg_partial_sum(reg_psum_17_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_12( .activation_in(reg_activation_17_11), .weight_in(reg_weight_16_12), .partial_sum_in(reg_psum_16_12), .reg_activation(reg_activation_17_12), .reg_weight(reg_weight_17_12), .reg_partial_sum(reg_psum_17_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_13( .activation_in(reg_activation_17_12), .weight_in(reg_weight_16_13), .partial_sum_in(reg_psum_16_13), .reg_activation(reg_activation_17_13), .reg_weight(reg_weight_17_13), .reg_partial_sum(reg_psum_17_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_14( .activation_in(reg_activation_17_13), .weight_in(reg_weight_16_14), .partial_sum_in(reg_psum_16_14), .reg_activation(reg_activation_17_14), .reg_weight(reg_weight_17_14), .reg_partial_sum(reg_psum_17_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_15( .activation_in(reg_activation_17_14), .weight_in(reg_weight_16_15), .partial_sum_in(reg_psum_16_15), .reg_activation(reg_activation_17_15), .reg_weight(reg_weight_17_15), .reg_partial_sum(reg_psum_17_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_16( .activation_in(reg_activation_17_15), .weight_in(reg_weight_16_16), .partial_sum_in(reg_psum_16_16), .reg_activation(reg_activation_17_16), .reg_weight(reg_weight_17_16), .reg_partial_sum(reg_psum_17_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_17( .activation_in(reg_activation_17_16), .weight_in(reg_weight_16_17), .partial_sum_in(reg_psum_16_17), .reg_activation(reg_activation_17_17), .reg_weight(reg_weight_17_17), .reg_partial_sum(reg_psum_17_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_18( .activation_in(reg_activation_17_17), .weight_in(reg_weight_16_18), .partial_sum_in(reg_psum_16_18), .reg_activation(reg_activation_17_18), .reg_weight(reg_weight_17_18), .reg_partial_sum(reg_psum_17_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_19( .activation_in(reg_activation_17_18), .weight_in(reg_weight_16_19), .partial_sum_in(reg_psum_16_19), .reg_activation(reg_activation_17_19), .reg_weight(reg_weight_17_19), .reg_partial_sum(reg_psum_17_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_20( .activation_in(reg_activation_17_19), .weight_in(reg_weight_16_20), .partial_sum_in(reg_psum_16_20), .reg_activation(reg_activation_17_20), .reg_weight(reg_weight_17_20), .reg_partial_sum(reg_psum_17_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_21( .activation_in(reg_activation_17_20), .weight_in(reg_weight_16_21), .partial_sum_in(reg_psum_16_21), .reg_activation(reg_activation_17_21), .reg_weight(reg_weight_17_21), .reg_partial_sum(reg_psum_17_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_22( .activation_in(reg_activation_17_21), .weight_in(reg_weight_16_22), .partial_sum_in(reg_psum_16_22), .reg_activation(reg_activation_17_22), .reg_weight(reg_weight_17_22), .reg_partial_sum(reg_psum_17_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_23( .activation_in(reg_activation_17_22), .weight_in(reg_weight_16_23), .partial_sum_in(reg_psum_16_23), .reg_activation(reg_activation_17_23), .reg_weight(reg_weight_17_23), .reg_partial_sum(reg_psum_17_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_24( .activation_in(reg_activation_17_23), .weight_in(reg_weight_16_24), .partial_sum_in(reg_psum_16_24), .reg_activation(reg_activation_17_24), .reg_weight(reg_weight_17_24), .reg_partial_sum(reg_psum_17_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_25( .activation_in(reg_activation_17_24), .weight_in(reg_weight_16_25), .partial_sum_in(reg_psum_16_25), .reg_activation(reg_activation_17_25), .reg_weight(reg_weight_17_25), .reg_partial_sum(reg_psum_17_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_26( .activation_in(reg_activation_17_25), .weight_in(reg_weight_16_26), .partial_sum_in(reg_psum_16_26), .reg_activation(reg_activation_17_26), .reg_weight(reg_weight_17_26), .reg_partial_sum(reg_psum_17_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_27( .activation_in(reg_activation_17_26), .weight_in(reg_weight_16_27), .partial_sum_in(reg_psum_16_27), .reg_activation(reg_activation_17_27), .reg_weight(reg_weight_17_27), .reg_partial_sum(reg_psum_17_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_28( .activation_in(reg_activation_17_27), .weight_in(reg_weight_16_28), .partial_sum_in(reg_psum_16_28), .reg_activation(reg_activation_17_28), .reg_weight(reg_weight_17_28), .reg_partial_sum(reg_psum_17_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_29( .activation_in(reg_activation_17_28), .weight_in(reg_weight_16_29), .partial_sum_in(reg_psum_16_29), .reg_activation(reg_activation_17_29), .reg_weight(reg_weight_17_29), .reg_partial_sum(reg_psum_17_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_30( .activation_in(reg_activation_17_29), .weight_in(reg_weight_16_30), .partial_sum_in(reg_psum_16_30), .reg_activation(reg_activation_17_30), .reg_weight(reg_weight_17_30), .reg_partial_sum(reg_psum_17_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_31( .activation_in(reg_activation_17_30), .weight_in(reg_weight_16_31), .partial_sum_in(reg_psum_16_31), .reg_activation(reg_activation_17_31), .reg_weight(reg_weight_17_31), .reg_partial_sum(reg_psum_17_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_32( .activation_in(reg_activation_17_31), .weight_in(reg_weight_16_32), .partial_sum_in(reg_psum_16_32), .reg_activation(reg_activation_17_32), .reg_weight(reg_weight_17_32), .reg_partial_sum(reg_psum_17_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_33( .activation_in(reg_activation_17_32), .weight_in(reg_weight_16_33), .partial_sum_in(reg_psum_16_33), .reg_activation(reg_activation_17_33), .reg_weight(reg_weight_17_33), .reg_partial_sum(reg_psum_17_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_34( .activation_in(reg_activation_17_33), .weight_in(reg_weight_16_34), .partial_sum_in(reg_psum_16_34), .reg_activation(reg_activation_17_34), .reg_weight(reg_weight_17_34), .reg_partial_sum(reg_psum_17_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_35( .activation_in(reg_activation_17_34), .weight_in(reg_weight_16_35), .partial_sum_in(reg_psum_16_35), .reg_activation(reg_activation_17_35), .reg_weight(reg_weight_17_35), .reg_partial_sum(reg_psum_17_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_36( .activation_in(reg_activation_17_35), .weight_in(reg_weight_16_36), .partial_sum_in(reg_psum_16_36), .reg_activation(reg_activation_17_36), .reg_weight(reg_weight_17_36), .reg_partial_sum(reg_psum_17_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_37( .activation_in(reg_activation_17_36), .weight_in(reg_weight_16_37), .partial_sum_in(reg_psum_16_37), .reg_activation(reg_activation_17_37), .reg_weight(reg_weight_17_37), .reg_partial_sum(reg_psum_17_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_38( .activation_in(reg_activation_17_37), .weight_in(reg_weight_16_38), .partial_sum_in(reg_psum_16_38), .reg_activation(reg_activation_17_38), .reg_weight(reg_weight_17_38), .reg_partial_sum(reg_psum_17_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_39( .activation_in(reg_activation_17_38), .weight_in(reg_weight_16_39), .partial_sum_in(reg_psum_16_39), .reg_activation(reg_activation_17_39), .reg_weight(reg_weight_17_39), .reg_partial_sum(reg_psum_17_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_40( .activation_in(reg_activation_17_39), .weight_in(reg_weight_16_40), .partial_sum_in(reg_psum_16_40), .reg_activation(reg_activation_17_40), .reg_weight(reg_weight_17_40), .reg_partial_sum(reg_psum_17_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_41( .activation_in(reg_activation_17_40), .weight_in(reg_weight_16_41), .partial_sum_in(reg_psum_16_41), .reg_activation(reg_activation_17_41), .reg_weight(reg_weight_17_41), .reg_partial_sum(reg_psum_17_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_42( .activation_in(reg_activation_17_41), .weight_in(reg_weight_16_42), .partial_sum_in(reg_psum_16_42), .reg_activation(reg_activation_17_42), .reg_weight(reg_weight_17_42), .reg_partial_sum(reg_psum_17_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_43( .activation_in(reg_activation_17_42), .weight_in(reg_weight_16_43), .partial_sum_in(reg_psum_16_43), .reg_activation(reg_activation_17_43), .reg_weight(reg_weight_17_43), .reg_partial_sum(reg_psum_17_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_44( .activation_in(reg_activation_17_43), .weight_in(reg_weight_16_44), .partial_sum_in(reg_psum_16_44), .reg_activation(reg_activation_17_44), .reg_weight(reg_weight_17_44), .reg_partial_sum(reg_psum_17_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_45( .activation_in(reg_activation_17_44), .weight_in(reg_weight_16_45), .partial_sum_in(reg_psum_16_45), .reg_activation(reg_activation_17_45), .reg_weight(reg_weight_17_45), .reg_partial_sum(reg_psum_17_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_46( .activation_in(reg_activation_17_45), .weight_in(reg_weight_16_46), .partial_sum_in(reg_psum_16_46), .reg_activation(reg_activation_17_46), .reg_weight(reg_weight_17_46), .reg_partial_sum(reg_psum_17_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_47( .activation_in(reg_activation_17_46), .weight_in(reg_weight_16_47), .partial_sum_in(reg_psum_16_47), .reg_activation(reg_activation_17_47), .reg_weight(reg_weight_17_47), .reg_partial_sum(reg_psum_17_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_48( .activation_in(reg_activation_17_47), .weight_in(reg_weight_16_48), .partial_sum_in(reg_psum_16_48), .reg_activation(reg_activation_17_48), .reg_weight(reg_weight_17_48), .reg_partial_sum(reg_psum_17_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_49( .activation_in(reg_activation_17_48), .weight_in(reg_weight_16_49), .partial_sum_in(reg_psum_16_49), .reg_activation(reg_activation_17_49), .reg_weight(reg_weight_17_49), .reg_partial_sum(reg_psum_17_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_50( .activation_in(reg_activation_17_49), .weight_in(reg_weight_16_50), .partial_sum_in(reg_psum_16_50), .reg_activation(reg_activation_17_50), .reg_weight(reg_weight_17_50), .reg_partial_sum(reg_psum_17_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_51( .activation_in(reg_activation_17_50), .weight_in(reg_weight_16_51), .partial_sum_in(reg_psum_16_51), .reg_activation(reg_activation_17_51), .reg_weight(reg_weight_17_51), .reg_partial_sum(reg_psum_17_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_52( .activation_in(reg_activation_17_51), .weight_in(reg_weight_16_52), .partial_sum_in(reg_psum_16_52), .reg_activation(reg_activation_17_52), .reg_weight(reg_weight_17_52), .reg_partial_sum(reg_psum_17_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_53( .activation_in(reg_activation_17_52), .weight_in(reg_weight_16_53), .partial_sum_in(reg_psum_16_53), .reg_activation(reg_activation_17_53), .reg_weight(reg_weight_17_53), .reg_partial_sum(reg_psum_17_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_54( .activation_in(reg_activation_17_53), .weight_in(reg_weight_16_54), .partial_sum_in(reg_psum_16_54), .reg_activation(reg_activation_17_54), .reg_weight(reg_weight_17_54), .reg_partial_sum(reg_psum_17_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_55( .activation_in(reg_activation_17_54), .weight_in(reg_weight_16_55), .partial_sum_in(reg_psum_16_55), .reg_activation(reg_activation_17_55), .reg_weight(reg_weight_17_55), .reg_partial_sum(reg_psum_17_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_56( .activation_in(reg_activation_17_55), .weight_in(reg_weight_16_56), .partial_sum_in(reg_psum_16_56), .reg_activation(reg_activation_17_56), .reg_weight(reg_weight_17_56), .reg_partial_sum(reg_psum_17_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_57( .activation_in(reg_activation_17_56), .weight_in(reg_weight_16_57), .partial_sum_in(reg_psum_16_57), .reg_activation(reg_activation_17_57), .reg_weight(reg_weight_17_57), .reg_partial_sum(reg_psum_17_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_58( .activation_in(reg_activation_17_57), .weight_in(reg_weight_16_58), .partial_sum_in(reg_psum_16_58), .reg_activation(reg_activation_17_58), .reg_weight(reg_weight_17_58), .reg_partial_sum(reg_psum_17_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_59( .activation_in(reg_activation_17_58), .weight_in(reg_weight_16_59), .partial_sum_in(reg_psum_16_59), .reg_activation(reg_activation_17_59), .reg_weight(reg_weight_17_59), .reg_partial_sum(reg_psum_17_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_60( .activation_in(reg_activation_17_59), .weight_in(reg_weight_16_60), .partial_sum_in(reg_psum_16_60), .reg_activation(reg_activation_17_60), .reg_weight(reg_weight_17_60), .reg_partial_sum(reg_psum_17_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_61( .activation_in(reg_activation_17_60), .weight_in(reg_weight_16_61), .partial_sum_in(reg_psum_16_61), .reg_activation(reg_activation_17_61), .reg_weight(reg_weight_17_61), .reg_partial_sum(reg_psum_17_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_62( .activation_in(reg_activation_17_61), .weight_in(reg_weight_16_62), .partial_sum_in(reg_psum_16_62), .reg_activation(reg_activation_17_62), .reg_weight(reg_weight_17_62), .reg_partial_sum(reg_psum_17_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_63( .activation_in(reg_activation_17_62), .weight_in(reg_weight_16_63), .partial_sum_in(reg_psum_16_63), .reg_weight(reg_weight_17_63), .reg_partial_sum(reg_psum_17_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_0( .activation_in(in_activation_18), .weight_in(reg_weight_17_0), .partial_sum_in(reg_psum_17_0), .reg_activation(reg_activation_18_0), .reg_weight(reg_weight_18_0), .reg_partial_sum(reg_psum_18_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_1( .activation_in(reg_activation_18_0), .weight_in(reg_weight_17_1), .partial_sum_in(reg_psum_17_1), .reg_activation(reg_activation_18_1), .reg_weight(reg_weight_18_1), .reg_partial_sum(reg_psum_18_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_2( .activation_in(reg_activation_18_1), .weight_in(reg_weight_17_2), .partial_sum_in(reg_psum_17_2), .reg_activation(reg_activation_18_2), .reg_weight(reg_weight_18_2), .reg_partial_sum(reg_psum_18_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_3( .activation_in(reg_activation_18_2), .weight_in(reg_weight_17_3), .partial_sum_in(reg_psum_17_3), .reg_activation(reg_activation_18_3), .reg_weight(reg_weight_18_3), .reg_partial_sum(reg_psum_18_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_4( .activation_in(reg_activation_18_3), .weight_in(reg_weight_17_4), .partial_sum_in(reg_psum_17_4), .reg_activation(reg_activation_18_4), .reg_weight(reg_weight_18_4), .reg_partial_sum(reg_psum_18_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_5( .activation_in(reg_activation_18_4), .weight_in(reg_weight_17_5), .partial_sum_in(reg_psum_17_5), .reg_activation(reg_activation_18_5), .reg_weight(reg_weight_18_5), .reg_partial_sum(reg_psum_18_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_6( .activation_in(reg_activation_18_5), .weight_in(reg_weight_17_6), .partial_sum_in(reg_psum_17_6), .reg_activation(reg_activation_18_6), .reg_weight(reg_weight_18_6), .reg_partial_sum(reg_psum_18_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_7( .activation_in(reg_activation_18_6), .weight_in(reg_weight_17_7), .partial_sum_in(reg_psum_17_7), .reg_activation(reg_activation_18_7), .reg_weight(reg_weight_18_7), .reg_partial_sum(reg_psum_18_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_8( .activation_in(reg_activation_18_7), .weight_in(reg_weight_17_8), .partial_sum_in(reg_psum_17_8), .reg_activation(reg_activation_18_8), .reg_weight(reg_weight_18_8), .reg_partial_sum(reg_psum_18_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_9( .activation_in(reg_activation_18_8), .weight_in(reg_weight_17_9), .partial_sum_in(reg_psum_17_9), .reg_activation(reg_activation_18_9), .reg_weight(reg_weight_18_9), .reg_partial_sum(reg_psum_18_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_10( .activation_in(reg_activation_18_9), .weight_in(reg_weight_17_10), .partial_sum_in(reg_psum_17_10), .reg_activation(reg_activation_18_10), .reg_weight(reg_weight_18_10), .reg_partial_sum(reg_psum_18_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_11( .activation_in(reg_activation_18_10), .weight_in(reg_weight_17_11), .partial_sum_in(reg_psum_17_11), .reg_activation(reg_activation_18_11), .reg_weight(reg_weight_18_11), .reg_partial_sum(reg_psum_18_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_12( .activation_in(reg_activation_18_11), .weight_in(reg_weight_17_12), .partial_sum_in(reg_psum_17_12), .reg_activation(reg_activation_18_12), .reg_weight(reg_weight_18_12), .reg_partial_sum(reg_psum_18_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_13( .activation_in(reg_activation_18_12), .weight_in(reg_weight_17_13), .partial_sum_in(reg_psum_17_13), .reg_activation(reg_activation_18_13), .reg_weight(reg_weight_18_13), .reg_partial_sum(reg_psum_18_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_14( .activation_in(reg_activation_18_13), .weight_in(reg_weight_17_14), .partial_sum_in(reg_psum_17_14), .reg_activation(reg_activation_18_14), .reg_weight(reg_weight_18_14), .reg_partial_sum(reg_psum_18_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_15( .activation_in(reg_activation_18_14), .weight_in(reg_weight_17_15), .partial_sum_in(reg_psum_17_15), .reg_activation(reg_activation_18_15), .reg_weight(reg_weight_18_15), .reg_partial_sum(reg_psum_18_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_16( .activation_in(reg_activation_18_15), .weight_in(reg_weight_17_16), .partial_sum_in(reg_psum_17_16), .reg_activation(reg_activation_18_16), .reg_weight(reg_weight_18_16), .reg_partial_sum(reg_psum_18_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_17( .activation_in(reg_activation_18_16), .weight_in(reg_weight_17_17), .partial_sum_in(reg_psum_17_17), .reg_activation(reg_activation_18_17), .reg_weight(reg_weight_18_17), .reg_partial_sum(reg_psum_18_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_18( .activation_in(reg_activation_18_17), .weight_in(reg_weight_17_18), .partial_sum_in(reg_psum_17_18), .reg_activation(reg_activation_18_18), .reg_weight(reg_weight_18_18), .reg_partial_sum(reg_psum_18_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_19( .activation_in(reg_activation_18_18), .weight_in(reg_weight_17_19), .partial_sum_in(reg_psum_17_19), .reg_activation(reg_activation_18_19), .reg_weight(reg_weight_18_19), .reg_partial_sum(reg_psum_18_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_20( .activation_in(reg_activation_18_19), .weight_in(reg_weight_17_20), .partial_sum_in(reg_psum_17_20), .reg_activation(reg_activation_18_20), .reg_weight(reg_weight_18_20), .reg_partial_sum(reg_psum_18_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_21( .activation_in(reg_activation_18_20), .weight_in(reg_weight_17_21), .partial_sum_in(reg_psum_17_21), .reg_activation(reg_activation_18_21), .reg_weight(reg_weight_18_21), .reg_partial_sum(reg_psum_18_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_22( .activation_in(reg_activation_18_21), .weight_in(reg_weight_17_22), .partial_sum_in(reg_psum_17_22), .reg_activation(reg_activation_18_22), .reg_weight(reg_weight_18_22), .reg_partial_sum(reg_psum_18_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_23( .activation_in(reg_activation_18_22), .weight_in(reg_weight_17_23), .partial_sum_in(reg_psum_17_23), .reg_activation(reg_activation_18_23), .reg_weight(reg_weight_18_23), .reg_partial_sum(reg_psum_18_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_24( .activation_in(reg_activation_18_23), .weight_in(reg_weight_17_24), .partial_sum_in(reg_psum_17_24), .reg_activation(reg_activation_18_24), .reg_weight(reg_weight_18_24), .reg_partial_sum(reg_psum_18_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_25( .activation_in(reg_activation_18_24), .weight_in(reg_weight_17_25), .partial_sum_in(reg_psum_17_25), .reg_activation(reg_activation_18_25), .reg_weight(reg_weight_18_25), .reg_partial_sum(reg_psum_18_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_26( .activation_in(reg_activation_18_25), .weight_in(reg_weight_17_26), .partial_sum_in(reg_psum_17_26), .reg_activation(reg_activation_18_26), .reg_weight(reg_weight_18_26), .reg_partial_sum(reg_psum_18_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_27( .activation_in(reg_activation_18_26), .weight_in(reg_weight_17_27), .partial_sum_in(reg_psum_17_27), .reg_activation(reg_activation_18_27), .reg_weight(reg_weight_18_27), .reg_partial_sum(reg_psum_18_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_28( .activation_in(reg_activation_18_27), .weight_in(reg_weight_17_28), .partial_sum_in(reg_psum_17_28), .reg_activation(reg_activation_18_28), .reg_weight(reg_weight_18_28), .reg_partial_sum(reg_psum_18_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_29( .activation_in(reg_activation_18_28), .weight_in(reg_weight_17_29), .partial_sum_in(reg_psum_17_29), .reg_activation(reg_activation_18_29), .reg_weight(reg_weight_18_29), .reg_partial_sum(reg_psum_18_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_30( .activation_in(reg_activation_18_29), .weight_in(reg_weight_17_30), .partial_sum_in(reg_psum_17_30), .reg_activation(reg_activation_18_30), .reg_weight(reg_weight_18_30), .reg_partial_sum(reg_psum_18_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_31( .activation_in(reg_activation_18_30), .weight_in(reg_weight_17_31), .partial_sum_in(reg_psum_17_31), .reg_activation(reg_activation_18_31), .reg_weight(reg_weight_18_31), .reg_partial_sum(reg_psum_18_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_32( .activation_in(reg_activation_18_31), .weight_in(reg_weight_17_32), .partial_sum_in(reg_psum_17_32), .reg_activation(reg_activation_18_32), .reg_weight(reg_weight_18_32), .reg_partial_sum(reg_psum_18_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_33( .activation_in(reg_activation_18_32), .weight_in(reg_weight_17_33), .partial_sum_in(reg_psum_17_33), .reg_activation(reg_activation_18_33), .reg_weight(reg_weight_18_33), .reg_partial_sum(reg_psum_18_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_34( .activation_in(reg_activation_18_33), .weight_in(reg_weight_17_34), .partial_sum_in(reg_psum_17_34), .reg_activation(reg_activation_18_34), .reg_weight(reg_weight_18_34), .reg_partial_sum(reg_psum_18_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_35( .activation_in(reg_activation_18_34), .weight_in(reg_weight_17_35), .partial_sum_in(reg_psum_17_35), .reg_activation(reg_activation_18_35), .reg_weight(reg_weight_18_35), .reg_partial_sum(reg_psum_18_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_36( .activation_in(reg_activation_18_35), .weight_in(reg_weight_17_36), .partial_sum_in(reg_psum_17_36), .reg_activation(reg_activation_18_36), .reg_weight(reg_weight_18_36), .reg_partial_sum(reg_psum_18_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_37( .activation_in(reg_activation_18_36), .weight_in(reg_weight_17_37), .partial_sum_in(reg_psum_17_37), .reg_activation(reg_activation_18_37), .reg_weight(reg_weight_18_37), .reg_partial_sum(reg_psum_18_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_38( .activation_in(reg_activation_18_37), .weight_in(reg_weight_17_38), .partial_sum_in(reg_psum_17_38), .reg_activation(reg_activation_18_38), .reg_weight(reg_weight_18_38), .reg_partial_sum(reg_psum_18_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_39( .activation_in(reg_activation_18_38), .weight_in(reg_weight_17_39), .partial_sum_in(reg_psum_17_39), .reg_activation(reg_activation_18_39), .reg_weight(reg_weight_18_39), .reg_partial_sum(reg_psum_18_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_40( .activation_in(reg_activation_18_39), .weight_in(reg_weight_17_40), .partial_sum_in(reg_psum_17_40), .reg_activation(reg_activation_18_40), .reg_weight(reg_weight_18_40), .reg_partial_sum(reg_psum_18_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_41( .activation_in(reg_activation_18_40), .weight_in(reg_weight_17_41), .partial_sum_in(reg_psum_17_41), .reg_activation(reg_activation_18_41), .reg_weight(reg_weight_18_41), .reg_partial_sum(reg_psum_18_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_42( .activation_in(reg_activation_18_41), .weight_in(reg_weight_17_42), .partial_sum_in(reg_psum_17_42), .reg_activation(reg_activation_18_42), .reg_weight(reg_weight_18_42), .reg_partial_sum(reg_psum_18_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_43( .activation_in(reg_activation_18_42), .weight_in(reg_weight_17_43), .partial_sum_in(reg_psum_17_43), .reg_activation(reg_activation_18_43), .reg_weight(reg_weight_18_43), .reg_partial_sum(reg_psum_18_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_44( .activation_in(reg_activation_18_43), .weight_in(reg_weight_17_44), .partial_sum_in(reg_psum_17_44), .reg_activation(reg_activation_18_44), .reg_weight(reg_weight_18_44), .reg_partial_sum(reg_psum_18_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_45( .activation_in(reg_activation_18_44), .weight_in(reg_weight_17_45), .partial_sum_in(reg_psum_17_45), .reg_activation(reg_activation_18_45), .reg_weight(reg_weight_18_45), .reg_partial_sum(reg_psum_18_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_46( .activation_in(reg_activation_18_45), .weight_in(reg_weight_17_46), .partial_sum_in(reg_psum_17_46), .reg_activation(reg_activation_18_46), .reg_weight(reg_weight_18_46), .reg_partial_sum(reg_psum_18_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_47( .activation_in(reg_activation_18_46), .weight_in(reg_weight_17_47), .partial_sum_in(reg_psum_17_47), .reg_activation(reg_activation_18_47), .reg_weight(reg_weight_18_47), .reg_partial_sum(reg_psum_18_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_48( .activation_in(reg_activation_18_47), .weight_in(reg_weight_17_48), .partial_sum_in(reg_psum_17_48), .reg_activation(reg_activation_18_48), .reg_weight(reg_weight_18_48), .reg_partial_sum(reg_psum_18_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_49( .activation_in(reg_activation_18_48), .weight_in(reg_weight_17_49), .partial_sum_in(reg_psum_17_49), .reg_activation(reg_activation_18_49), .reg_weight(reg_weight_18_49), .reg_partial_sum(reg_psum_18_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_50( .activation_in(reg_activation_18_49), .weight_in(reg_weight_17_50), .partial_sum_in(reg_psum_17_50), .reg_activation(reg_activation_18_50), .reg_weight(reg_weight_18_50), .reg_partial_sum(reg_psum_18_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_51( .activation_in(reg_activation_18_50), .weight_in(reg_weight_17_51), .partial_sum_in(reg_psum_17_51), .reg_activation(reg_activation_18_51), .reg_weight(reg_weight_18_51), .reg_partial_sum(reg_psum_18_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_52( .activation_in(reg_activation_18_51), .weight_in(reg_weight_17_52), .partial_sum_in(reg_psum_17_52), .reg_activation(reg_activation_18_52), .reg_weight(reg_weight_18_52), .reg_partial_sum(reg_psum_18_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_53( .activation_in(reg_activation_18_52), .weight_in(reg_weight_17_53), .partial_sum_in(reg_psum_17_53), .reg_activation(reg_activation_18_53), .reg_weight(reg_weight_18_53), .reg_partial_sum(reg_psum_18_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_54( .activation_in(reg_activation_18_53), .weight_in(reg_weight_17_54), .partial_sum_in(reg_psum_17_54), .reg_activation(reg_activation_18_54), .reg_weight(reg_weight_18_54), .reg_partial_sum(reg_psum_18_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_55( .activation_in(reg_activation_18_54), .weight_in(reg_weight_17_55), .partial_sum_in(reg_psum_17_55), .reg_activation(reg_activation_18_55), .reg_weight(reg_weight_18_55), .reg_partial_sum(reg_psum_18_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_56( .activation_in(reg_activation_18_55), .weight_in(reg_weight_17_56), .partial_sum_in(reg_psum_17_56), .reg_activation(reg_activation_18_56), .reg_weight(reg_weight_18_56), .reg_partial_sum(reg_psum_18_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_57( .activation_in(reg_activation_18_56), .weight_in(reg_weight_17_57), .partial_sum_in(reg_psum_17_57), .reg_activation(reg_activation_18_57), .reg_weight(reg_weight_18_57), .reg_partial_sum(reg_psum_18_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_58( .activation_in(reg_activation_18_57), .weight_in(reg_weight_17_58), .partial_sum_in(reg_psum_17_58), .reg_activation(reg_activation_18_58), .reg_weight(reg_weight_18_58), .reg_partial_sum(reg_psum_18_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_59( .activation_in(reg_activation_18_58), .weight_in(reg_weight_17_59), .partial_sum_in(reg_psum_17_59), .reg_activation(reg_activation_18_59), .reg_weight(reg_weight_18_59), .reg_partial_sum(reg_psum_18_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_60( .activation_in(reg_activation_18_59), .weight_in(reg_weight_17_60), .partial_sum_in(reg_psum_17_60), .reg_activation(reg_activation_18_60), .reg_weight(reg_weight_18_60), .reg_partial_sum(reg_psum_18_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_61( .activation_in(reg_activation_18_60), .weight_in(reg_weight_17_61), .partial_sum_in(reg_psum_17_61), .reg_activation(reg_activation_18_61), .reg_weight(reg_weight_18_61), .reg_partial_sum(reg_psum_18_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_62( .activation_in(reg_activation_18_61), .weight_in(reg_weight_17_62), .partial_sum_in(reg_psum_17_62), .reg_activation(reg_activation_18_62), .reg_weight(reg_weight_18_62), .reg_partial_sum(reg_psum_18_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_63( .activation_in(reg_activation_18_62), .weight_in(reg_weight_17_63), .partial_sum_in(reg_psum_17_63), .reg_weight(reg_weight_18_63), .reg_partial_sum(reg_psum_18_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_0( .activation_in(in_activation_19), .weight_in(reg_weight_18_0), .partial_sum_in(reg_psum_18_0), .reg_activation(reg_activation_19_0), .reg_weight(reg_weight_19_0), .reg_partial_sum(reg_psum_19_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_1( .activation_in(reg_activation_19_0), .weight_in(reg_weight_18_1), .partial_sum_in(reg_psum_18_1), .reg_activation(reg_activation_19_1), .reg_weight(reg_weight_19_1), .reg_partial_sum(reg_psum_19_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_2( .activation_in(reg_activation_19_1), .weight_in(reg_weight_18_2), .partial_sum_in(reg_psum_18_2), .reg_activation(reg_activation_19_2), .reg_weight(reg_weight_19_2), .reg_partial_sum(reg_psum_19_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_3( .activation_in(reg_activation_19_2), .weight_in(reg_weight_18_3), .partial_sum_in(reg_psum_18_3), .reg_activation(reg_activation_19_3), .reg_weight(reg_weight_19_3), .reg_partial_sum(reg_psum_19_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_4( .activation_in(reg_activation_19_3), .weight_in(reg_weight_18_4), .partial_sum_in(reg_psum_18_4), .reg_activation(reg_activation_19_4), .reg_weight(reg_weight_19_4), .reg_partial_sum(reg_psum_19_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_5( .activation_in(reg_activation_19_4), .weight_in(reg_weight_18_5), .partial_sum_in(reg_psum_18_5), .reg_activation(reg_activation_19_5), .reg_weight(reg_weight_19_5), .reg_partial_sum(reg_psum_19_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_6( .activation_in(reg_activation_19_5), .weight_in(reg_weight_18_6), .partial_sum_in(reg_psum_18_6), .reg_activation(reg_activation_19_6), .reg_weight(reg_weight_19_6), .reg_partial_sum(reg_psum_19_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_7( .activation_in(reg_activation_19_6), .weight_in(reg_weight_18_7), .partial_sum_in(reg_psum_18_7), .reg_activation(reg_activation_19_7), .reg_weight(reg_weight_19_7), .reg_partial_sum(reg_psum_19_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_8( .activation_in(reg_activation_19_7), .weight_in(reg_weight_18_8), .partial_sum_in(reg_psum_18_8), .reg_activation(reg_activation_19_8), .reg_weight(reg_weight_19_8), .reg_partial_sum(reg_psum_19_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_9( .activation_in(reg_activation_19_8), .weight_in(reg_weight_18_9), .partial_sum_in(reg_psum_18_9), .reg_activation(reg_activation_19_9), .reg_weight(reg_weight_19_9), .reg_partial_sum(reg_psum_19_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_10( .activation_in(reg_activation_19_9), .weight_in(reg_weight_18_10), .partial_sum_in(reg_psum_18_10), .reg_activation(reg_activation_19_10), .reg_weight(reg_weight_19_10), .reg_partial_sum(reg_psum_19_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_11( .activation_in(reg_activation_19_10), .weight_in(reg_weight_18_11), .partial_sum_in(reg_psum_18_11), .reg_activation(reg_activation_19_11), .reg_weight(reg_weight_19_11), .reg_partial_sum(reg_psum_19_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_12( .activation_in(reg_activation_19_11), .weight_in(reg_weight_18_12), .partial_sum_in(reg_psum_18_12), .reg_activation(reg_activation_19_12), .reg_weight(reg_weight_19_12), .reg_partial_sum(reg_psum_19_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_13( .activation_in(reg_activation_19_12), .weight_in(reg_weight_18_13), .partial_sum_in(reg_psum_18_13), .reg_activation(reg_activation_19_13), .reg_weight(reg_weight_19_13), .reg_partial_sum(reg_psum_19_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_14( .activation_in(reg_activation_19_13), .weight_in(reg_weight_18_14), .partial_sum_in(reg_psum_18_14), .reg_activation(reg_activation_19_14), .reg_weight(reg_weight_19_14), .reg_partial_sum(reg_psum_19_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_15( .activation_in(reg_activation_19_14), .weight_in(reg_weight_18_15), .partial_sum_in(reg_psum_18_15), .reg_activation(reg_activation_19_15), .reg_weight(reg_weight_19_15), .reg_partial_sum(reg_psum_19_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_16( .activation_in(reg_activation_19_15), .weight_in(reg_weight_18_16), .partial_sum_in(reg_psum_18_16), .reg_activation(reg_activation_19_16), .reg_weight(reg_weight_19_16), .reg_partial_sum(reg_psum_19_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_17( .activation_in(reg_activation_19_16), .weight_in(reg_weight_18_17), .partial_sum_in(reg_psum_18_17), .reg_activation(reg_activation_19_17), .reg_weight(reg_weight_19_17), .reg_partial_sum(reg_psum_19_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_18( .activation_in(reg_activation_19_17), .weight_in(reg_weight_18_18), .partial_sum_in(reg_psum_18_18), .reg_activation(reg_activation_19_18), .reg_weight(reg_weight_19_18), .reg_partial_sum(reg_psum_19_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_19( .activation_in(reg_activation_19_18), .weight_in(reg_weight_18_19), .partial_sum_in(reg_psum_18_19), .reg_activation(reg_activation_19_19), .reg_weight(reg_weight_19_19), .reg_partial_sum(reg_psum_19_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_20( .activation_in(reg_activation_19_19), .weight_in(reg_weight_18_20), .partial_sum_in(reg_psum_18_20), .reg_activation(reg_activation_19_20), .reg_weight(reg_weight_19_20), .reg_partial_sum(reg_psum_19_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_21( .activation_in(reg_activation_19_20), .weight_in(reg_weight_18_21), .partial_sum_in(reg_psum_18_21), .reg_activation(reg_activation_19_21), .reg_weight(reg_weight_19_21), .reg_partial_sum(reg_psum_19_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_22( .activation_in(reg_activation_19_21), .weight_in(reg_weight_18_22), .partial_sum_in(reg_psum_18_22), .reg_activation(reg_activation_19_22), .reg_weight(reg_weight_19_22), .reg_partial_sum(reg_psum_19_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_23( .activation_in(reg_activation_19_22), .weight_in(reg_weight_18_23), .partial_sum_in(reg_psum_18_23), .reg_activation(reg_activation_19_23), .reg_weight(reg_weight_19_23), .reg_partial_sum(reg_psum_19_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_24( .activation_in(reg_activation_19_23), .weight_in(reg_weight_18_24), .partial_sum_in(reg_psum_18_24), .reg_activation(reg_activation_19_24), .reg_weight(reg_weight_19_24), .reg_partial_sum(reg_psum_19_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_25( .activation_in(reg_activation_19_24), .weight_in(reg_weight_18_25), .partial_sum_in(reg_psum_18_25), .reg_activation(reg_activation_19_25), .reg_weight(reg_weight_19_25), .reg_partial_sum(reg_psum_19_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_26( .activation_in(reg_activation_19_25), .weight_in(reg_weight_18_26), .partial_sum_in(reg_psum_18_26), .reg_activation(reg_activation_19_26), .reg_weight(reg_weight_19_26), .reg_partial_sum(reg_psum_19_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_27( .activation_in(reg_activation_19_26), .weight_in(reg_weight_18_27), .partial_sum_in(reg_psum_18_27), .reg_activation(reg_activation_19_27), .reg_weight(reg_weight_19_27), .reg_partial_sum(reg_psum_19_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_28( .activation_in(reg_activation_19_27), .weight_in(reg_weight_18_28), .partial_sum_in(reg_psum_18_28), .reg_activation(reg_activation_19_28), .reg_weight(reg_weight_19_28), .reg_partial_sum(reg_psum_19_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_29( .activation_in(reg_activation_19_28), .weight_in(reg_weight_18_29), .partial_sum_in(reg_psum_18_29), .reg_activation(reg_activation_19_29), .reg_weight(reg_weight_19_29), .reg_partial_sum(reg_psum_19_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_30( .activation_in(reg_activation_19_29), .weight_in(reg_weight_18_30), .partial_sum_in(reg_psum_18_30), .reg_activation(reg_activation_19_30), .reg_weight(reg_weight_19_30), .reg_partial_sum(reg_psum_19_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_31( .activation_in(reg_activation_19_30), .weight_in(reg_weight_18_31), .partial_sum_in(reg_psum_18_31), .reg_activation(reg_activation_19_31), .reg_weight(reg_weight_19_31), .reg_partial_sum(reg_psum_19_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_32( .activation_in(reg_activation_19_31), .weight_in(reg_weight_18_32), .partial_sum_in(reg_psum_18_32), .reg_activation(reg_activation_19_32), .reg_weight(reg_weight_19_32), .reg_partial_sum(reg_psum_19_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_33( .activation_in(reg_activation_19_32), .weight_in(reg_weight_18_33), .partial_sum_in(reg_psum_18_33), .reg_activation(reg_activation_19_33), .reg_weight(reg_weight_19_33), .reg_partial_sum(reg_psum_19_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_34( .activation_in(reg_activation_19_33), .weight_in(reg_weight_18_34), .partial_sum_in(reg_psum_18_34), .reg_activation(reg_activation_19_34), .reg_weight(reg_weight_19_34), .reg_partial_sum(reg_psum_19_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_35( .activation_in(reg_activation_19_34), .weight_in(reg_weight_18_35), .partial_sum_in(reg_psum_18_35), .reg_activation(reg_activation_19_35), .reg_weight(reg_weight_19_35), .reg_partial_sum(reg_psum_19_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_36( .activation_in(reg_activation_19_35), .weight_in(reg_weight_18_36), .partial_sum_in(reg_psum_18_36), .reg_activation(reg_activation_19_36), .reg_weight(reg_weight_19_36), .reg_partial_sum(reg_psum_19_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_37( .activation_in(reg_activation_19_36), .weight_in(reg_weight_18_37), .partial_sum_in(reg_psum_18_37), .reg_activation(reg_activation_19_37), .reg_weight(reg_weight_19_37), .reg_partial_sum(reg_psum_19_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_38( .activation_in(reg_activation_19_37), .weight_in(reg_weight_18_38), .partial_sum_in(reg_psum_18_38), .reg_activation(reg_activation_19_38), .reg_weight(reg_weight_19_38), .reg_partial_sum(reg_psum_19_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_39( .activation_in(reg_activation_19_38), .weight_in(reg_weight_18_39), .partial_sum_in(reg_psum_18_39), .reg_activation(reg_activation_19_39), .reg_weight(reg_weight_19_39), .reg_partial_sum(reg_psum_19_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_40( .activation_in(reg_activation_19_39), .weight_in(reg_weight_18_40), .partial_sum_in(reg_psum_18_40), .reg_activation(reg_activation_19_40), .reg_weight(reg_weight_19_40), .reg_partial_sum(reg_psum_19_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_41( .activation_in(reg_activation_19_40), .weight_in(reg_weight_18_41), .partial_sum_in(reg_psum_18_41), .reg_activation(reg_activation_19_41), .reg_weight(reg_weight_19_41), .reg_partial_sum(reg_psum_19_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_42( .activation_in(reg_activation_19_41), .weight_in(reg_weight_18_42), .partial_sum_in(reg_psum_18_42), .reg_activation(reg_activation_19_42), .reg_weight(reg_weight_19_42), .reg_partial_sum(reg_psum_19_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_43( .activation_in(reg_activation_19_42), .weight_in(reg_weight_18_43), .partial_sum_in(reg_psum_18_43), .reg_activation(reg_activation_19_43), .reg_weight(reg_weight_19_43), .reg_partial_sum(reg_psum_19_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_44( .activation_in(reg_activation_19_43), .weight_in(reg_weight_18_44), .partial_sum_in(reg_psum_18_44), .reg_activation(reg_activation_19_44), .reg_weight(reg_weight_19_44), .reg_partial_sum(reg_psum_19_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_45( .activation_in(reg_activation_19_44), .weight_in(reg_weight_18_45), .partial_sum_in(reg_psum_18_45), .reg_activation(reg_activation_19_45), .reg_weight(reg_weight_19_45), .reg_partial_sum(reg_psum_19_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_46( .activation_in(reg_activation_19_45), .weight_in(reg_weight_18_46), .partial_sum_in(reg_psum_18_46), .reg_activation(reg_activation_19_46), .reg_weight(reg_weight_19_46), .reg_partial_sum(reg_psum_19_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_47( .activation_in(reg_activation_19_46), .weight_in(reg_weight_18_47), .partial_sum_in(reg_psum_18_47), .reg_activation(reg_activation_19_47), .reg_weight(reg_weight_19_47), .reg_partial_sum(reg_psum_19_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_48( .activation_in(reg_activation_19_47), .weight_in(reg_weight_18_48), .partial_sum_in(reg_psum_18_48), .reg_activation(reg_activation_19_48), .reg_weight(reg_weight_19_48), .reg_partial_sum(reg_psum_19_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_49( .activation_in(reg_activation_19_48), .weight_in(reg_weight_18_49), .partial_sum_in(reg_psum_18_49), .reg_activation(reg_activation_19_49), .reg_weight(reg_weight_19_49), .reg_partial_sum(reg_psum_19_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_50( .activation_in(reg_activation_19_49), .weight_in(reg_weight_18_50), .partial_sum_in(reg_psum_18_50), .reg_activation(reg_activation_19_50), .reg_weight(reg_weight_19_50), .reg_partial_sum(reg_psum_19_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_51( .activation_in(reg_activation_19_50), .weight_in(reg_weight_18_51), .partial_sum_in(reg_psum_18_51), .reg_activation(reg_activation_19_51), .reg_weight(reg_weight_19_51), .reg_partial_sum(reg_psum_19_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_52( .activation_in(reg_activation_19_51), .weight_in(reg_weight_18_52), .partial_sum_in(reg_psum_18_52), .reg_activation(reg_activation_19_52), .reg_weight(reg_weight_19_52), .reg_partial_sum(reg_psum_19_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_53( .activation_in(reg_activation_19_52), .weight_in(reg_weight_18_53), .partial_sum_in(reg_psum_18_53), .reg_activation(reg_activation_19_53), .reg_weight(reg_weight_19_53), .reg_partial_sum(reg_psum_19_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_54( .activation_in(reg_activation_19_53), .weight_in(reg_weight_18_54), .partial_sum_in(reg_psum_18_54), .reg_activation(reg_activation_19_54), .reg_weight(reg_weight_19_54), .reg_partial_sum(reg_psum_19_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_55( .activation_in(reg_activation_19_54), .weight_in(reg_weight_18_55), .partial_sum_in(reg_psum_18_55), .reg_activation(reg_activation_19_55), .reg_weight(reg_weight_19_55), .reg_partial_sum(reg_psum_19_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_56( .activation_in(reg_activation_19_55), .weight_in(reg_weight_18_56), .partial_sum_in(reg_psum_18_56), .reg_activation(reg_activation_19_56), .reg_weight(reg_weight_19_56), .reg_partial_sum(reg_psum_19_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_57( .activation_in(reg_activation_19_56), .weight_in(reg_weight_18_57), .partial_sum_in(reg_psum_18_57), .reg_activation(reg_activation_19_57), .reg_weight(reg_weight_19_57), .reg_partial_sum(reg_psum_19_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_58( .activation_in(reg_activation_19_57), .weight_in(reg_weight_18_58), .partial_sum_in(reg_psum_18_58), .reg_activation(reg_activation_19_58), .reg_weight(reg_weight_19_58), .reg_partial_sum(reg_psum_19_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_59( .activation_in(reg_activation_19_58), .weight_in(reg_weight_18_59), .partial_sum_in(reg_psum_18_59), .reg_activation(reg_activation_19_59), .reg_weight(reg_weight_19_59), .reg_partial_sum(reg_psum_19_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_60( .activation_in(reg_activation_19_59), .weight_in(reg_weight_18_60), .partial_sum_in(reg_psum_18_60), .reg_activation(reg_activation_19_60), .reg_weight(reg_weight_19_60), .reg_partial_sum(reg_psum_19_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_61( .activation_in(reg_activation_19_60), .weight_in(reg_weight_18_61), .partial_sum_in(reg_psum_18_61), .reg_activation(reg_activation_19_61), .reg_weight(reg_weight_19_61), .reg_partial_sum(reg_psum_19_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_62( .activation_in(reg_activation_19_61), .weight_in(reg_weight_18_62), .partial_sum_in(reg_psum_18_62), .reg_activation(reg_activation_19_62), .reg_weight(reg_weight_19_62), .reg_partial_sum(reg_psum_19_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_63( .activation_in(reg_activation_19_62), .weight_in(reg_weight_18_63), .partial_sum_in(reg_psum_18_63), .reg_weight(reg_weight_19_63), .reg_partial_sum(reg_psum_19_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_0( .activation_in(in_activation_20), .weight_in(reg_weight_19_0), .partial_sum_in(reg_psum_19_0), .reg_activation(reg_activation_20_0), .reg_weight(reg_weight_20_0), .reg_partial_sum(reg_psum_20_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_1( .activation_in(reg_activation_20_0), .weight_in(reg_weight_19_1), .partial_sum_in(reg_psum_19_1), .reg_activation(reg_activation_20_1), .reg_weight(reg_weight_20_1), .reg_partial_sum(reg_psum_20_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_2( .activation_in(reg_activation_20_1), .weight_in(reg_weight_19_2), .partial_sum_in(reg_psum_19_2), .reg_activation(reg_activation_20_2), .reg_weight(reg_weight_20_2), .reg_partial_sum(reg_psum_20_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_3( .activation_in(reg_activation_20_2), .weight_in(reg_weight_19_3), .partial_sum_in(reg_psum_19_3), .reg_activation(reg_activation_20_3), .reg_weight(reg_weight_20_3), .reg_partial_sum(reg_psum_20_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_4( .activation_in(reg_activation_20_3), .weight_in(reg_weight_19_4), .partial_sum_in(reg_psum_19_4), .reg_activation(reg_activation_20_4), .reg_weight(reg_weight_20_4), .reg_partial_sum(reg_psum_20_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_5( .activation_in(reg_activation_20_4), .weight_in(reg_weight_19_5), .partial_sum_in(reg_psum_19_5), .reg_activation(reg_activation_20_5), .reg_weight(reg_weight_20_5), .reg_partial_sum(reg_psum_20_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_6( .activation_in(reg_activation_20_5), .weight_in(reg_weight_19_6), .partial_sum_in(reg_psum_19_6), .reg_activation(reg_activation_20_6), .reg_weight(reg_weight_20_6), .reg_partial_sum(reg_psum_20_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_7( .activation_in(reg_activation_20_6), .weight_in(reg_weight_19_7), .partial_sum_in(reg_psum_19_7), .reg_activation(reg_activation_20_7), .reg_weight(reg_weight_20_7), .reg_partial_sum(reg_psum_20_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_8( .activation_in(reg_activation_20_7), .weight_in(reg_weight_19_8), .partial_sum_in(reg_psum_19_8), .reg_activation(reg_activation_20_8), .reg_weight(reg_weight_20_8), .reg_partial_sum(reg_psum_20_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_9( .activation_in(reg_activation_20_8), .weight_in(reg_weight_19_9), .partial_sum_in(reg_psum_19_9), .reg_activation(reg_activation_20_9), .reg_weight(reg_weight_20_9), .reg_partial_sum(reg_psum_20_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_10( .activation_in(reg_activation_20_9), .weight_in(reg_weight_19_10), .partial_sum_in(reg_psum_19_10), .reg_activation(reg_activation_20_10), .reg_weight(reg_weight_20_10), .reg_partial_sum(reg_psum_20_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_11( .activation_in(reg_activation_20_10), .weight_in(reg_weight_19_11), .partial_sum_in(reg_psum_19_11), .reg_activation(reg_activation_20_11), .reg_weight(reg_weight_20_11), .reg_partial_sum(reg_psum_20_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_12( .activation_in(reg_activation_20_11), .weight_in(reg_weight_19_12), .partial_sum_in(reg_psum_19_12), .reg_activation(reg_activation_20_12), .reg_weight(reg_weight_20_12), .reg_partial_sum(reg_psum_20_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_13( .activation_in(reg_activation_20_12), .weight_in(reg_weight_19_13), .partial_sum_in(reg_psum_19_13), .reg_activation(reg_activation_20_13), .reg_weight(reg_weight_20_13), .reg_partial_sum(reg_psum_20_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_14( .activation_in(reg_activation_20_13), .weight_in(reg_weight_19_14), .partial_sum_in(reg_psum_19_14), .reg_activation(reg_activation_20_14), .reg_weight(reg_weight_20_14), .reg_partial_sum(reg_psum_20_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_15( .activation_in(reg_activation_20_14), .weight_in(reg_weight_19_15), .partial_sum_in(reg_psum_19_15), .reg_activation(reg_activation_20_15), .reg_weight(reg_weight_20_15), .reg_partial_sum(reg_psum_20_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_16( .activation_in(reg_activation_20_15), .weight_in(reg_weight_19_16), .partial_sum_in(reg_psum_19_16), .reg_activation(reg_activation_20_16), .reg_weight(reg_weight_20_16), .reg_partial_sum(reg_psum_20_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_17( .activation_in(reg_activation_20_16), .weight_in(reg_weight_19_17), .partial_sum_in(reg_psum_19_17), .reg_activation(reg_activation_20_17), .reg_weight(reg_weight_20_17), .reg_partial_sum(reg_psum_20_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_18( .activation_in(reg_activation_20_17), .weight_in(reg_weight_19_18), .partial_sum_in(reg_psum_19_18), .reg_activation(reg_activation_20_18), .reg_weight(reg_weight_20_18), .reg_partial_sum(reg_psum_20_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_19( .activation_in(reg_activation_20_18), .weight_in(reg_weight_19_19), .partial_sum_in(reg_psum_19_19), .reg_activation(reg_activation_20_19), .reg_weight(reg_weight_20_19), .reg_partial_sum(reg_psum_20_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_20( .activation_in(reg_activation_20_19), .weight_in(reg_weight_19_20), .partial_sum_in(reg_psum_19_20), .reg_activation(reg_activation_20_20), .reg_weight(reg_weight_20_20), .reg_partial_sum(reg_psum_20_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_21( .activation_in(reg_activation_20_20), .weight_in(reg_weight_19_21), .partial_sum_in(reg_psum_19_21), .reg_activation(reg_activation_20_21), .reg_weight(reg_weight_20_21), .reg_partial_sum(reg_psum_20_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_22( .activation_in(reg_activation_20_21), .weight_in(reg_weight_19_22), .partial_sum_in(reg_psum_19_22), .reg_activation(reg_activation_20_22), .reg_weight(reg_weight_20_22), .reg_partial_sum(reg_psum_20_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_23( .activation_in(reg_activation_20_22), .weight_in(reg_weight_19_23), .partial_sum_in(reg_psum_19_23), .reg_activation(reg_activation_20_23), .reg_weight(reg_weight_20_23), .reg_partial_sum(reg_psum_20_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_24( .activation_in(reg_activation_20_23), .weight_in(reg_weight_19_24), .partial_sum_in(reg_psum_19_24), .reg_activation(reg_activation_20_24), .reg_weight(reg_weight_20_24), .reg_partial_sum(reg_psum_20_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_25( .activation_in(reg_activation_20_24), .weight_in(reg_weight_19_25), .partial_sum_in(reg_psum_19_25), .reg_activation(reg_activation_20_25), .reg_weight(reg_weight_20_25), .reg_partial_sum(reg_psum_20_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_26( .activation_in(reg_activation_20_25), .weight_in(reg_weight_19_26), .partial_sum_in(reg_psum_19_26), .reg_activation(reg_activation_20_26), .reg_weight(reg_weight_20_26), .reg_partial_sum(reg_psum_20_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_27( .activation_in(reg_activation_20_26), .weight_in(reg_weight_19_27), .partial_sum_in(reg_psum_19_27), .reg_activation(reg_activation_20_27), .reg_weight(reg_weight_20_27), .reg_partial_sum(reg_psum_20_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_28( .activation_in(reg_activation_20_27), .weight_in(reg_weight_19_28), .partial_sum_in(reg_psum_19_28), .reg_activation(reg_activation_20_28), .reg_weight(reg_weight_20_28), .reg_partial_sum(reg_psum_20_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_29( .activation_in(reg_activation_20_28), .weight_in(reg_weight_19_29), .partial_sum_in(reg_psum_19_29), .reg_activation(reg_activation_20_29), .reg_weight(reg_weight_20_29), .reg_partial_sum(reg_psum_20_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_30( .activation_in(reg_activation_20_29), .weight_in(reg_weight_19_30), .partial_sum_in(reg_psum_19_30), .reg_activation(reg_activation_20_30), .reg_weight(reg_weight_20_30), .reg_partial_sum(reg_psum_20_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_31( .activation_in(reg_activation_20_30), .weight_in(reg_weight_19_31), .partial_sum_in(reg_psum_19_31), .reg_activation(reg_activation_20_31), .reg_weight(reg_weight_20_31), .reg_partial_sum(reg_psum_20_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_32( .activation_in(reg_activation_20_31), .weight_in(reg_weight_19_32), .partial_sum_in(reg_psum_19_32), .reg_activation(reg_activation_20_32), .reg_weight(reg_weight_20_32), .reg_partial_sum(reg_psum_20_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_33( .activation_in(reg_activation_20_32), .weight_in(reg_weight_19_33), .partial_sum_in(reg_psum_19_33), .reg_activation(reg_activation_20_33), .reg_weight(reg_weight_20_33), .reg_partial_sum(reg_psum_20_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_34( .activation_in(reg_activation_20_33), .weight_in(reg_weight_19_34), .partial_sum_in(reg_psum_19_34), .reg_activation(reg_activation_20_34), .reg_weight(reg_weight_20_34), .reg_partial_sum(reg_psum_20_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_35( .activation_in(reg_activation_20_34), .weight_in(reg_weight_19_35), .partial_sum_in(reg_psum_19_35), .reg_activation(reg_activation_20_35), .reg_weight(reg_weight_20_35), .reg_partial_sum(reg_psum_20_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_36( .activation_in(reg_activation_20_35), .weight_in(reg_weight_19_36), .partial_sum_in(reg_psum_19_36), .reg_activation(reg_activation_20_36), .reg_weight(reg_weight_20_36), .reg_partial_sum(reg_psum_20_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_37( .activation_in(reg_activation_20_36), .weight_in(reg_weight_19_37), .partial_sum_in(reg_psum_19_37), .reg_activation(reg_activation_20_37), .reg_weight(reg_weight_20_37), .reg_partial_sum(reg_psum_20_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_38( .activation_in(reg_activation_20_37), .weight_in(reg_weight_19_38), .partial_sum_in(reg_psum_19_38), .reg_activation(reg_activation_20_38), .reg_weight(reg_weight_20_38), .reg_partial_sum(reg_psum_20_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_39( .activation_in(reg_activation_20_38), .weight_in(reg_weight_19_39), .partial_sum_in(reg_psum_19_39), .reg_activation(reg_activation_20_39), .reg_weight(reg_weight_20_39), .reg_partial_sum(reg_psum_20_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_40( .activation_in(reg_activation_20_39), .weight_in(reg_weight_19_40), .partial_sum_in(reg_psum_19_40), .reg_activation(reg_activation_20_40), .reg_weight(reg_weight_20_40), .reg_partial_sum(reg_psum_20_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_41( .activation_in(reg_activation_20_40), .weight_in(reg_weight_19_41), .partial_sum_in(reg_psum_19_41), .reg_activation(reg_activation_20_41), .reg_weight(reg_weight_20_41), .reg_partial_sum(reg_psum_20_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_42( .activation_in(reg_activation_20_41), .weight_in(reg_weight_19_42), .partial_sum_in(reg_psum_19_42), .reg_activation(reg_activation_20_42), .reg_weight(reg_weight_20_42), .reg_partial_sum(reg_psum_20_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_43( .activation_in(reg_activation_20_42), .weight_in(reg_weight_19_43), .partial_sum_in(reg_psum_19_43), .reg_activation(reg_activation_20_43), .reg_weight(reg_weight_20_43), .reg_partial_sum(reg_psum_20_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_44( .activation_in(reg_activation_20_43), .weight_in(reg_weight_19_44), .partial_sum_in(reg_psum_19_44), .reg_activation(reg_activation_20_44), .reg_weight(reg_weight_20_44), .reg_partial_sum(reg_psum_20_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_45( .activation_in(reg_activation_20_44), .weight_in(reg_weight_19_45), .partial_sum_in(reg_psum_19_45), .reg_activation(reg_activation_20_45), .reg_weight(reg_weight_20_45), .reg_partial_sum(reg_psum_20_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_46( .activation_in(reg_activation_20_45), .weight_in(reg_weight_19_46), .partial_sum_in(reg_psum_19_46), .reg_activation(reg_activation_20_46), .reg_weight(reg_weight_20_46), .reg_partial_sum(reg_psum_20_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_47( .activation_in(reg_activation_20_46), .weight_in(reg_weight_19_47), .partial_sum_in(reg_psum_19_47), .reg_activation(reg_activation_20_47), .reg_weight(reg_weight_20_47), .reg_partial_sum(reg_psum_20_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_48( .activation_in(reg_activation_20_47), .weight_in(reg_weight_19_48), .partial_sum_in(reg_psum_19_48), .reg_activation(reg_activation_20_48), .reg_weight(reg_weight_20_48), .reg_partial_sum(reg_psum_20_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_49( .activation_in(reg_activation_20_48), .weight_in(reg_weight_19_49), .partial_sum_in(reg_psum_19_49), .reg_activation(reg_activation_20_49), .reg_weight(reg_weight_20_49), .reg_partial_sum(reg_psum_20_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_50( .activation_in(reg_activation_20_49), .weight_in(reg_weight_19_50), .partial_sum_in(reg_psum_19_50), .reg_activation(reg_activation_20_50), .reg_weight(reg_weight_20_50), .reg_partial_sum(reg_psum_20_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_51( .activation_in(reg_activation_20_50), .weight_in(reg_weight_19_51), .partial_sum_in(reg_psum_19_51), .reg_activation(reg_activation_20_51), .reg_weight(reg_weight_20_51), .reg_partial_sum(reg_psum_20_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_52( .activation_in(reg_activation_20_51), .weight_in(reg_weight_19_52), .partial_sum_in(reg_psum_19_52), .reg_activation(reg_activation_20_52), .reg_weight(reg_weight_20_52), .reg_partial_sum(reg_psum_20_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_53( .activation_in(reg_activation_20_52), .weight_in(reg_weight_19_53), .partial_sum_in(reg_psum_19_53), .reg_activation(reg_activation_20_53), .reg_weight(reg_weight_20_53), .reg_partial_sum(reg_psum_20_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_54( .activation_in(reg_activation_20_53), .weight_in(reg_weight_19_54), .partial_sum_in(reg_psum_19_54), .reg_activation(reg_activation_20_54), .reg_weight(reg_weight_20_54), .reg_partial_sum(reg_psum_20_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_55( .activation_in(reg_activation_20_54), .weight_in(reg_weight_19_55), .partial_sum_in(reg_psum_19_55), .reg_activation(reg_activation_20_55), .reg_weight(reg_weight_20_55), .reg_partial_sum(reg_psum_20_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_56( .activation_in(reg_activation_20_55), .weight_in(reg_weight_19_56), .partial_sum_in(reg_psum_19_56), .reg_activation(reg_activation_20_56), .reg_weight(reg_weight_20_56), .reg_partial_sum(reg_psum_20_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_57( .activation_in(reg_activation_20_56), .weight_in(reg_weight_19_57), .partial_sum_in(reg_psum_19_57), .reg_activation(reg_activation_20_57), .reg_weight(reg_weight_20_57), .reg_partial_sum(reg_psum_20_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_58( .activation_in(reg_activation_20_57), .weight_in(reg_weight_19_58), .partial_sum_in(reg_psum_19_58), .reg_activation(reg_activation_20_58), .reg_weight(reg_weight_20_58), .reg_partial_sum(reg_psum_20_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_59( .activation_in(reg_activation_20_58), .weight_in(reg_weight_19_59), .partial_sum_in(reg_psum_19_59), .reg_activation(reg_activation_20_59), .reg_weight(reg_weight_20_59), .reg_partial_sum(reg_psum_20_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_60( .activation_in(reg_activation_20_59), .weight_in(reg_weight_19_60), .partial_sum_in(reg_psum_19_60), .reg_activation(reg_activation_20_60), .reg_weight(reg_weight_20_60), .reg_partial_sum(reg_psum_20_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_61( .activation_in(reg_activation_20_60), .weight_in(reg_weight_19_61), .partial_sum_in(reg_psum_19_61), .reg_activation(reg_activation_20_61), .reg_weight(reg_weight_20_61), .reg_partial_sum(reg_psum_20_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_62( .activation_in(reg_activation_20_61), .weight_in(reg_weight_19_62), .partial_sum_in(reg_psum_19_62), .reg_activation(reg_activation_20_62), .reg_weight(reg_weight_20_62), .reg_partial_sum(reg_psum_20_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_63( .activation_in(reg_activation_20_62), .weight_in(reg_weight_19_63), .partial_sum_in(reg_psum_19_63), .reg_weight(reg_weight_20_63), .reg_partial_sum(reg_psum_20_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_0( .activation_in(in_activation_21), .weight_in(reg_weight_20_0), .partial_sum_in(reg_psum_20_0), .reg_activation(reg_activation_21_0), .reg_weight(reg_weight_21_0), .reg_partial_sum(reg_psum_21_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_1( .activation_in(reg_activation_21_0), .weight_in(reg_weight_20_1), .partial_sum_in(reg_psum_20_1), .reg_activation(reg_activation_21_1), .reg_weight(reg_weight_21_1), .reg_partial_sum(reg_psum_21_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_2( .activation_in(reg_activation_21_1), .weight_in(reg_weight_20_2), .partial_sum_in(reg_psum_20_2), .reg_activation(reg_activation_21_2), .reg_weight(reg_weight_21_2), .reg_partial_sum(reg_psum_21_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_3( .activation_in(reg_activation_21_2), .weight_in(reg_weight_20_3), .partial_sum_in(reg_psum_20_3), .reg_activation(reg_activation_21_3), .reg_weight(reg_weight_21_3), .reg_partial_sum(reg_psum_21_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_4( .activation_in(reg_activation_21_3), .weight_in(reg_weight_20_4), .partial_sum_in(reg_psum_20_4), .reg_activation(reg_activation_21_4), .reg_weight(reg_weight_21_4), .reg_partial_sum(reg_psum_21_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_5( .activation_in(reg_activation_21_4), .weight_in(reg_weight_20_5), .partial_sum_in(reg_psum_20_5), .reg_activation(reg_activation_21_5), .reg_weight(reg_weight_21_5), .reg_partial_sum(reg_psum_21_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_6( .activation_in(reg_activation_21_5), .weight_in(reg_weight_20_6), .partial_sum_in(reg_psum_20_6), .reg_activation(reg_activation_21_6), .reg_weight(reg_weight_21_6), .reg_partial_sum(reg_psum_21_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_7( .activation_in(reg_activation_21_6), .weight_in(reg_weight_20_7), .partial_sum_in(reg_psum_20_7), .reg_activation(reg_activation_21_7), .reg_weight(reg_weight_21_7), .reg_partial_sum(reg_psum_21_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_8( .activation_in(reg_activation_21_7), .weight_in(reg_weight_20_8), .partial_sum_in(reg_psum_20_8), .reg_activation(reg_activation_21_8), .reg_weight(reg_weight_21_8), .reg_partial_sum(reg_psum_21_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_9( .activation_in(reg_activation_21_8), .weight_in(reg_weight_20_9), .partial_sum_in(reg_psum_20_9), .reg_activation(reg_activation_21_9), .reg_weight(reg_weight_21_9), .reg_partial_sum(reg_psum_21_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_10( .activation_in(reg_activation_21_9), .weight_in(reg_weight_20_10), .partial_sum_in(reg_psum_20_10), .reg_activation(reg_activation_21_10), .reg_weight(reg_weight_21_10), .reg_partial_sum(reg_psum_21_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_11( .activation_in(reg_activation_21_10), .weight_in(reg_weight_20_11), .partial_sum_in(reg_psum_20_11), .reg_activation(reg_activation_21_11), .reg_weight(reg_weight_21_11), .reg_partial_sum(reg_psum_21_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_12( .activation_in(reg_activation_21_11), .weight_in(reg_weight_20_12), .partial_sum_in(reg_psum_20_12), .reg_activation(reg_activation_21_12), .reg_weight(reg_weight_21_12), .reg_partial_sum(reg_psum_21_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_13( .activation_in(reg_activation_21_12), .weight_in(reg_weight_20_13), .partial_sum_in(reg_psum_20_13), .reg_activation(reg_activation_21_13), .reg_weight(reg_weight_21_13), .reg_partial_sum(reg_psum_21_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_14( .activation_in(reg_activation_21_13), .weight_in(reg_weight_20_14), .partial_sum_in(reg_psum_20_14), .reg_activation(reg_activation_21_14), .reg_weight(reg_weight_21_14), .reg_partial_sum(reg_psum_21_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_15( .activation_in(reg_activation_21_14), .weight_in(reg_weight_20_15), .partial_sum_in(reg_psum_20_15), .reg_activation(reg_activation_21_15), .reg_weight(reg_weight_21_15), .reg_partial_sum(reg_psum_21_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_16( .activation_in(reg_activation_21_15), .weight_in(reg_weight_20_16), .partial_sum_in(reg_psum_20_16), .reg_activation(reg_activation_21_16), .reg_weight(reg_weight_21_16), .reg_partial_sum(reg_psum_21_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_17( .activation_in(reg_activation_21_16), .weight_in(reg_weight_20_17), .partial_sum_in(reg_psum_20_17), .reg_activation(reg_activation_21_17), .reg_weight(reg_weight_21_17), .reg_partial_sum(reg_psum_21_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_18( .activation_in(reg_activation_21_17), .weight_in(reg_weight_20_18), .partial_sum_in(reg_psum_20_18), .reg_activation(reg_activation_21_18), .reg_weight(reg_weight_21_18), .reg_partial_sum(reg_psum_21_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_19( .activation_in(reg_activation_21_18), .weight_in(reg_weight_20_19), .partial_sum_in(reg_psum_20_19), .reg_activation(reg_activation_21_19), .reg_weight(reg_weight_21_19), .reg_partial_sum(reg_psum_21_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_20( .activation_in(reg_activation_21_19), .weight_in(reg_weight_20_20), .partial_sum_in(reg_psum_20_20), .reg_activation(reg_activation_21_20), .reg_weight(reg_weight_21_20), .reg_partial_sum(reg_psum_21_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_21( .activation_in(reg_activation_21_20), .weight_in(reg_weight_20_21), .partial_sum_in(reg_psum_20_21), .reg_activation(reg_activation_21_21), .reg_weight(reg_weight_21_21), .reg_partial_sum(reg_psum_21_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_22( .activation_in(reg_activation_21_21), .weight_in(reg_weight_20_22), .partial_sum_in(reg_psum_20_22), .reg_activation(reg_activation_21_22), .reg_weight(reg_weight_21_22), .reg_partial_sum(reg_psum_21_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_23( .activation_in(reg_activation_21_22), .weight_in(reg_weight_20_23), .partial_sum_in(reg_psum_20_23), .reg_activation(reg_activation_21_23), .reg_weight(reg_weight_21_23), .reg_partial_sum(reg_psum_21_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_24( .activation_in(reg_activation_21_23), .weight_in(reg_weight_20_24), .partial_sum_in(reg_psum_20_24), .reg_activation(reg_activation_21_24), .reg_weight(reg_weight_21_24), .reg_partial_sum(reg_psum_21_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_25( .activation_in(reg_activation_21_24), .weight_in(reg_weight_20_25), .partial_sum_in(reg_psum_20_25), .reg_activation(reg_activation_21_25), .reg_weight(reg_weight_21_25), .reg_partial_sum(reg_psum_21_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_26( .activation_in(reg_activation_21_25), .weight_in(reg_weight_20_26), .partial_sum_in(reg_psum_20_26), .reg_activation(reg_activation_21_26), .reg_weight(reg_weight_21_26), .reg_partial_sum(reg_psum_21_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_27( .activation_in(reg_activation_21_26), .weight_in(reg_weight_20_27), .partial_sum_in(reg_psum_20_27), .reg_activation(reg_activation_21_27), .reg_weight(reg_weight_21_27), .reg_partial_sum(reg_psum_21_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_28( .activation_in(reg_activation_21_27), .weight_in(reg_weight_20_28), .partial_sum_in(reg_psum_20_28), .reg_activation(reg_activation_21_28), .reg_weight(reg_weight_21_28), .reg_partial_sum(reg_psum_21_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_29( .activation_in(reg_activation_21_28), .weight_in(reg_weight_20_29), .partial_sum_in(reg_psum_20_29), .reg_activation(reg_activation_21_29), .reg_weight(reg_weight_21_29), .reg_partial_sum(reg_psum_21_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_30( .activation_in(reg_activation_21_29), .weight_in(reg_weight_20_30), .partial_sum_in(reg_psum_20_30), .reg_activation(reg_activation_21_30), .reg_weight(reg_weight_21_30), .reg_partial_sum(reg_psum_21_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_31( .activation_in(reg_activation_21_30), .weight_in(reg_weight_20_31), .partial_sum_in(reg_psum_20_31), .reg_activation(reg_activation_21_31), .reg_weight(reg_weight_21_31), .reg_partial_sum(reg_psum_21_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_32( .activation_in(reg_activation_21_31), .weight_in(reg_weight_20_32), .partial_sum_in(reg_psum_20_32), .reg_activation(reg_activation_21_32), .reg_weight(reg_weight_21_32), .reg_partial_sum(reg_psum_21_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_33( .activation_in(reg_activation_21_32), .weight_in(reg_weight_20_33), .partial_sum_in(reg_psum_20_33), .reg_activation(reg_activation_21_33), .reg_weight(reg_weight_21_33), .reg_partial_sum(reg_psum_21_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_34( .activation_in(reg_activation_21_33), .weight_in(reg_weight_20_34), .partial_sum_in(reg_psum_20_34), .reg_activation(reg_activation_21_34), .reg_weight(reg_weight_21_34), .reg_partial_sum(reg_psum_21_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_35( .activation_in(reg_activation_21_34), .weight_in(reg_weight_20_35), .partial_sum_in(reg_psum_20_35), .reg_activation(reg_activation_21_35), .reg_weight(reg_weight_21_35), .reg_partial_sum(reg_psum_21_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_36( .activation_in(reg_activation_21_35), .weight_in(reg_weight_20_36), .partial_sum_in(reg_psum_20_36), .reg_activation(reg_activation_21_36), .reg_weight(reg_weight_21_36), .reg_partial_sum(reg_psum_21_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_37( .activation_in(reg_activation_21_36), .weight_in(reg_weight_20_37), .partial_sum_in(reg_psum_20_37), .reg_activation(reg_activation_21_37), .reg_weight(reg_weight_21_37), .reg_partial_sum(reg_psum_21_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_38( .activation_in(reg_activation_21_37), .weight_in(reg_weight_20_38), .partial_sum_in(reg_psum_20_38), .reg_activation(reg_activation_21_38), .reg_weight(reg_weight_21_38), .reg_partial_sum(reg_psum_21_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_39( .activation_in(reg_activation_21_38), .weight_in(reg_weight_20_39), .partial_sum_in(reg_psum_20_39), .reg_activation(reg_activation_21_39), .reg_weight(reg_weight_21_39), .reg_partial_sum(reg_psum_21_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_40( .activation_in(reg_activation_21_39), .weight_in(reg_weight_20_40), .partial_sum_in(reg_psum_20_40), .reg_activation(reg_activation_21_40), .reg_weight(reg_weight_21_40), .reg_partial_sum(reg_psum_21_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_41( .activation_in(reg_activation_21_40), .weight_in(reg_weight_20_41), .partial_sum_in(reg_psum_20_41), .reg_activation(reg_activation_21_41), .reg_weight(reg_weight_21_41), .reg_partial_sum(reg_psum_21_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_42( .activation_in(reg_activation_21_41), .weight_in(reg_weight_20_42), .partial_sum_in(reg_psum_20_42), .reg_activation(reg_activation_21_42), .reg_weight(reg_weight_21_42), .reg_partial_sum(reg_psum_21_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_43( .activation_in(reg_activation_21_42), .weight_in(reg_weight_20_43), .partial_sum_in(reg_psum_20_43), .reg_activation(reg_activation_21_43), .reg_weight(reg_weight_21_43), .reg_partial_sum(reg_psum_21_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_44( .activation_in(reg_activation_21_43), .weight_in(reg_weight_20_44), .partial_sum_in(reg_psum_20_44), .reg_activation(reg_activation_21_44), .reg_weight(reg_weight_21_44), .reg_partial_sum(reg_psum_21_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_45( .activation_in(reg_activation_21_44), .weight_in(reg_weight_20_45), .partial_sum_in(reg_psum_20_45), .reg_activation(reg_activation_21_45), .reg_weight(reg_weight_21_45), .reg_partial_sum(reg_psum_21_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_46( .activation_in(reg_activation_21_45), .weight_in(reg_weight_20_46), .partial_sum_in(reg_psum_20_46), .reg_activation(reg_activation_21_46), .reg_weight(reg_weight_21_46), .reg_partial_sum(reg_psum_21_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_47( .activation_in(reg_activation_21_46), .weight_in(reg_weight_20_47), .partial_sum_in(reg_psum_20_47), .reg_activation(reg_activation_21_47), .reg_weight(reg_weight_21_47), .reg_partial_sum(reg_psum_21_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_48( .activation_in(reg_activation_21_47), .weight_in(reg_weight_20_48), .partial_sum_in(reg_psum_20_48), .reg_activation(reg_activation_21_48), .reg_weight(reg_weight_21_48), .reg_partial_sum(reg_psum_21_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_49( .activation_in(reg_activation_21_48), .weight_in(reg_weight_20_49), .partial_sum_in(reg_psum_20_49), .reg_activation(reg_activation_21_49), .reg_weight(reg_weight_21_49), .reg_partial_sum(reg_psum_21_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_50( .activation_in(reg_activation_21_49), .weight_in(reg_weight_20_50), .partial_sum_in(reg_psum_20_50), .reg_activation(reg_activation_21_50), .reg_weight(reg_weight_21_50), .reg_partial_sum(reg_psum_21_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_51( .activation_in(reg_activation_21_50), .weight_in(reg_weight_20_51), .partial_sum_in(reg_psum_20_51), .reg_activation(reg_activation_21_51), .reg_weight(reg_weight_21_51), .reg_partial_sum(reg_psum_21_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_52( .activation_in(reg_activation_21_51), .weight_in(reg_weight_20_52), .partial_sum_in(reg_psum_20_52), .reg_activation(reg_activation_21_52), .reg_weight(reg_weight_21_52), .reg_partial_sum(reg_psum_21_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_53( .activation_in(reg_activation_21_52), .weight_in(reg_weight_20_53), .partial_sum_in(reg_psum_20_53), .reg_activation(reg_activation_21_53), .reg_weight(reg_weight_21_53), .reg_partial_sum(reg_psum_21_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_54( .activation_in(reg_activation_21_53), .weight_in(reg_weight_20_54), .partial_sum_in(reg_psum_20_54), .reg_activation(reg_activation_21_54), .reg_weight(reg_weight_21_54), .reg_partial_sum(reg_psum_21_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_55( .activation_in(reg_activation_21_54), .weight_in(reg_weight_20_55), .partial_sum_in(reg_psum_20_55), .reg_activation(reg_activation_21_55), .reg_weight(reg_weight_21_55), .reg_partial_sum(reg_psum_21_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_56( .activation_in(reg_activation_21_55), .weight_in(reg_weight_20_56), .partial_sum_in(reg_psum_20_56), .reg_activation(reg_activation_21_56), .reg_weight(reg_weight_21_56), .reg_partial_sum(reg_psum_21_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_57( .activation_in(reg_activation_21_56), .weight_in(reg_weight_20_57), .partial_sum_in(reg_psum_20_57), .reg_activation(reg_activation_21_57), .reg_weight(reg_weight_21_57), .reg_partial_sum(reg_psum_21_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_58( .activation_in(reg_activation_21_57), .weight_in(reg_weight_20_58), .partial_sum_in(reg_psum_20_58), .reg_activation(reg_activation_21_58), .reg_weight(reg_weight_21_58), .reg_partial_sum(reg_psum_21_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_59( .activation_in(reg_activation_21_58), .weight_in(reg_weight_20_59), .partial_sum_in(reg_psum_20_59), .reg_activation(reg_activation_21_59), .reg_weight(reg_weight_21_59), .reg_partial_sum(reg_psum_21_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_60( .activation_in(reg_activation_21_59), .weight_in(reg_weight_20_60), .partial_sum_in(reg_psum_20_60), .reg_activation(reg_activation_21_60), .reg_weight(reg_weight_21_60), .reg_partial_sum(reg_psum_21_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_61( .activation_in(reg_activation_21_60), .weight_in(reg_weight_20_61), .partial_sum_in(reg_psum_20_61), .reg_activation(reg_activation_21_61), .reg_weight(reg_weight_21_61), .reg_partial_sum(reg_psum_21_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_62( .activation_in(reg_activation_21_61), .weight_in(reg_weight_20_62), .partial_sum_in(reg_psum_20_62), .reg_activation(reg_activation_21_62), .reg_weight(reg_weight_21_62), .reg_partial_sum(reg_psum_21_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_63( .activation_in(reg_activation_21_62), .weight_in(reg_weight_20_63), .partial_sum_in(reg_psum_20_63), .reg_weight(reg_weight_21_63), .reg_partial_sum(reg_psum_21_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_0( .activation_in(in_activation_22), .weight_in(reg_weight_21_0), .partial_sum_in(reg_psum_21_0), .reg_activation(reg_activation_22_0), .reg_weight(reg_weight_22_0), .reg_partial_sum(reg_psum_22_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_1( .activation_in(reg_activation_22_0), .weight_in(reg_weight_21_1), .partial_sum_in(reg_psum_21_1), .reg_activation(reg_activation_22_1), .reg_weight(reg_weight_22_1), .reg_partial_sum(reg_psum_22_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_2( .activation_in(reg_activation_22_1), .weight_in(reg_weight_21_2), .partial_sum_in(reg_psum_21_2), .reg_activation(reg_activation_22_2), .reg_weight(reg_weight_22_2), .reg_partial_sum(reg_psum_22_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_3( .activation_in(reg_activation_22_2), .weight_in(reg_weight_21_3), .partial_sum_in(reg_psum_21_3), .reg_activation(reg_activation_22_3), .reg_weight(reg_weight_22_3), .reg_partial_sum(reg_psum_22_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_4( .activation_in(reg_activation_22_3), .weight_in(reg_weight_21_4), .partial_sum_in(reg_psum_21_4), .reg_activation(reg_activation_22_4), .reg_weight(reg_weight_22_4), .reg_partial_sum(reg_psum_22_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_5( .activation_in(reg_activation_22_4), .weight_in(reg_weight_21_5), .partial_sum_in(reg_psum_21_5), .reg_activation(reg_activation_22_5), .reg_weight(reg_weight_22_5), .reg_partial_sum(reg_psum_22_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_6( .activation_in(reg_activation_22_5), .weight_in(reg_weight_21_6), .partial_sum_in(reg_psum_21_6), .reg_activation(reg_activation_22_6), .reg_weight(reg_weight_22_6), .reg_partial_sum(reg_psum_22_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_7( .activation_in(reg_activation_22_6), .weight_in(reg_weight_21_7), .partial_sum_in(reg_psum_21_7), .reg_activation(reg_activation_22_7), .reg_weight(reg_weight_22_7), .reg_partial_sum(reg_psum_22_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_8( .activation_in(reg_activation_22_7), .weight_in(reg_weight_21_8), .partial_sum_in(reg_psum_21_8), .reg_activation(reg_activation_22_8), .reg_weight(reg_weight_22_8), .reg_partial_sum(reg_psum_22_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_9( .activation_in(reg_activation_22_8), .weight_in(reg_weight_21_9), .partial_sum_in(reg_psum_21_9), .reg_activation(reg_activation_22_9), .reg_weight(reg_weight_22_9), .reg_partial_sum(reg_psum_22_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_10( .activation_in(reg_activation_22_9), .weight_in(reg_weight_21_10), .partial_sum_in(reg_psum_21_10), .reg_activation(reg_activation_22_10), .reg_weight(reg_weight_22_10), .reg_partial_sum(reg_psum_22_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_11( .activation_in(reg_activation_22_10), .weight_in(reg_weight_21_11), .partial_sum_in(reg_psum_21_11), .reg_activation(reg_activation_22_11), .reg_weight(reg_weight_22_11), .reg_partial_sum(reg_psum_22_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_12( .activation_in(reg_activation_22_11), .weight_in(reg_weight_21_12), .partial_sum_in(reg_psum_21_12), .reg_activation(reg_activation_22_12), .reg_weight(reg_weight_22_12), .reg_partial_sum(reg_psum_22_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_13( .activation_in(reg_activation_22_12), .weight_in(reg_weight_21_13), .partial_sum_in(reg_psum_21_13), .reg_activation(reg_activation_22_13), .reg_weight(reg_weight_22_13), .reg_partial_sum(reg_psum_22_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_14( .activation_in(reg_activation_22_13), .weight_in(reg_weight_21_14), .partial_sum_in(reg_psum_21_14), .reg_activation(reg_activation_22_14), .reg_weight(reg_weight_22_14), .reg_partial_sum(reg_psum_22_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_15( .activation_in(reg_activation_22_14), .weight_in(reg_weight_21_15), .partial_sum_in(reg_psum_21_15), .reg_activation(reg_activation_22_15), .reg_weight(reg_weight_22_15), .reg_partial_sum(reg_psum_22_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_16( .activation_in(reg_activation_22_15), .weight_in(reg_weight_21_16), .partial_sum_in(reg_psum_21_16), .reg_activation(reg_activation_22_16), .reg_weight(reg_weight_22_16), .reg_partial_sum(reg_psum_22_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_17( .activation_in(reg_activation_22_16), .weight_in(reg_weight_21_17), .partial_sum_in(reg_psum_21_17), .reg_activation(reg_activation_22_17), .reg_weight(reg_weight_22_17), .reg_partial_sum(reg_psum_22_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_18( .activation_in(reg_activation_22_17), .weight_in(reg_weight_21_18), .partial_sum_in(reg_psum_21_18), .reg_activation(reg_activation_22_18), .reg_weight(reg_weight_22_18), .reg_partial_sum(reg_psum_22_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_19( .activation_in(reg_activation_22_18), .weight_in(reg_weight_21_19), .partial_sum_in(reg_psum_21_19), .reg_activation(reg_activation_22_19), .reg_weight(reg_weight_22_19), .reg_partial_sum(reg_psum_22_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_20( .activation_in(reg_activation_22_19), .weight_in(reg_weight_21_20), .partial_sum_in(reg_psum_21_20), .reg_activation(reg_activation_22_20), .reg_weight(reg_weight_22_20), .reg_partial_sum(reg_psum_22_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_21( .activation_in(reg_activation_22_20), .weight_in(reg_weight_21_21), .partial_sum_in(reg_psum_21_21), .reg_activation(reg_activation_22_21), .reg_weight(reg_weight_22_21), .reg_partial_sum(reg_psum_22_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_22( .activation_in(reg_activation_22_21), .weight_in(reg_weight_21_22), .partial_sum_in(reg_psum_21_22), .reg_activation(reg_activation_22_22), .reg_weight(reg_weight_22_22), .reg_partial_sum(reg_psum_22_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_23( .activation_in(reg_activation_22_22), .weight_in(reg_weight_21_23), .partial_sum_in(reg_psum_21_23), .reg_activation(reg_activation_22_23), .reg_weight(reg_weight_22_23), .reg_partial_sum(reg_psum_22_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_24( .activation_in(reg_activation_22_23), .weight_in(reg_weight_21_24), .partial_sum_in(reg_psum_21_24), .reg_activation(reg_activation_22_24), .reg_weight(reg_weight_22_24), .reg_partial_sum(reg_psum_22_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_25( .activation_in(reg_activation_22_24), .weight_in(reg_weight_21_25), .partial_sum_in(reg_psum_21_25), .reg_activation(reg_activation_22_25), .reg_weight(reg_weight_22_25), .reg_partial_sum(reg_psum_22_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_26( .activation_in(reg_activation_22_25), .weight_in(reg_weight_21_26), .partial_sum_in(reg_psum_21_26), .reg_activation(reg_activation_22_26), .reg_weight(reg_weight_22_26), .reg_partial_sum(reg_psum_22_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_27( .activation_in(reg_activation_22_26), .weight_in(reg_weight_21_27), .partial_sum_in(reg_psum_21_27), .reg_activation(reg_activation_22_27), .reg_weight(reg_weight_22_27), .reg_partial_sum(reg_psum_22_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_28( .activation_in(reg_activation_22_27), .weight_in(reg_weight_21_28), .partial_sum_in(reg_psum_21_28), .reg_activation(reg_activation_22_28), .reg_weight(reg_weight_22_28), .reg_partial_sum(reg_psum_22_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_29( .activation_in(reg_activation_22_28), .weight_in(reg_weight_21_29), .partial_sum_in(reg_psum_21_29), .reg_activation(reg_activation_22_29), .reg_weight(reg_weight_22_29), .reg_partial_sum(reg_psum_22_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_30( .activation_in(reg_activation_22_29), .weight_in(reg_weight_21_30), .partial_sum_in(reg_psum_21_30), .reg_activation(reg_activation_22_30), .reg_weight(reg_weight_22_30), .reg_partial_sum(reg_psum_22_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_31( .activation_in(reg_activation_22_30), .weight_in(reg_weight_21_31), .partial_sum_in(reg_psum_21_31), .reg_activation(reg_activation_22_31), .reg_weight(reg_weight_22_31), .reg_partial_sum(reg_psum_22_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_32( .activation_in(reg_activation_22_31), .weight_in(reg_weight_21_32), .partial_sum_in(reg_psum_21_32), .reg_activation(reg_activation_22_32), .reg_weight(reg_weight_22_32), .reg_partial_sum(reg_psum_22_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_33( .activation_in(reg_activation_22_32), .weight_in(reg_weight_21_33), .partial_sum_in(reg_psum_21_33), .reg_activation(reg_activation_22_33), .reg_weight(reg_weight_22_33), .reg_partial_sum(reg_psum_22_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_34( .activation_in(reg_activation_22_33), .weight_in(reg_weight_21_34), .partial_sum_in(reg_psum_21_34), .reg_activation(reg_activation_22_34), .reg_weight(reg_weight_22_34), .reg_partial_sum(reg_psum_22_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_35( .activation_in(reg_activation_22_34), .weight_in(reg_weight_21_35), .partial_sum_in(reg_psum_21_35), .reg_activation(reg_activation_22_35), .reg_weight(reg_weight_22_35), .reg_partial_sum(reg_psum_22_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_36( .activation_in(reg_activation_22_35), .weight_in(reg_weight_21_36), .partial_sum_in(reg_psum_21_36), .reg_activation(reg_activation_22_36), .reg_weight(reg_weight_22_36), .reg_partial_sum(reg_psum_22_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_37( .activation_in(reg_activation_22_36), .weight_in(reg_weight_21_37), .partial_sum_in(reg_psum_21_37), .reg_activation(reg_activation_22_37), .reg_weight(reg_weight_22_37), .reg_partial_sum(reg_psum_22_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_38( .activation_in(reg_activation_22_37), .weight_in(reg_weight_21_38), .partial_sum_in(reg_psum_21_38), .reg_activation(reg_activation_22_38), .reg_weight(reg_weight_22_38), .reg_partial_sum(reg_psum_22_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_39( .activation_in(reg_activation_22_38), .weight_in(reg_weight_21_39), .partial_sum_in(reg_psum_21_39), .reg_activation(reg_activation_22_39), .reg_weight(reg_weight_22_39), .reg_partial_sum(reg_psum_22_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_40( .activation_in(reg_activation_22_39), .weight_in(reg_weight_21_40), .partial_sum_in(reg_psum_21_40), .reg_activation(reg_activation_22_40), .reg_weight(reg_weight_22_40), .reg_partial_sum(reg_psum_22_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_41( .activation_in(reg_activation_22_40), .weight_in(reg_weight_21_41), .partial_sum_in(reg_psum_21_41), .reg_activation(reg_activation_22_41), .reg_weight(reg_weight_22_41), .reg_partial_sum(reg_psum_22_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_42( .activation_in(reg_activation_22_41), .weight_in(reg_weight_21_42), .partial_sum_in(reg_psum_21_42), .reg_activation(reg_activation_22_42), .reg_weight(reg_weight_22_42), .reg_partial_sum(reg_psum_22_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_43( .activation_in(reg_activation_22_42), .weight_in(reg_weight_21_43), .partial_sum_in(reg_psum_21_43), .reg_activation(reg_activation_22_43), .reg_weight(reg_weight_22_43), .reg_partial_sum(reg_psum_22_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_44( .activation_in(reg_activation_22_43), .weight_in(reg_weight_21_44), .partial_sum_in(reg_psum_21_44), .reg_activation(reg_activation_22_44), .reg_weight(reg_weight_22_44), .reg_partial_sum(reg_psum_22_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_45( .activation_in(reg_activation_22_44), .weight_in(reg_weight_21_45), .partial_sum_in(reg_psum_21_45), .reg_activation(reg_activation_22_45), .reg_weight(reg_weight_22_45), .reg_partial_sum(reg_psum_22_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_46( .activation_in(reg_activation_22_45), .weight_in(reg_weight_21_46), .partial_sum_in(reg_psum_21_46), .reg_activation(reg_activation_22_46), .reg_weight(reg_weight_22_46), .reg_partial_sum(reg_psum_22_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_47( .activation_in(reg_activation_22_46), .weight_in(reg_weight_21_47), .partial_sum_in(reg_psum_21_47), .reg_activation(reg_activation_22_47), .reg_weight(reg_weight_22_47), .reg_partial_sum(reg_psum_22_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_48( .activation_in(reg_activation_22_47), .weight_in(reg_weight_21_48), .partial_sum_in(reg_psum_21_48), .reg_activation(reg_activation_22_48), .reg_weight(reg_weight_22_48), .reg_partial_sum(reg_psum_22_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_49( .activation_in(reg_activation_22_48), .weight_in(reg_weight_21_49), .partial_sum_in(reg_psum_21_49), .reg_activation(reg_activation_22_49), .reg_weight(reg_weight_22_49), .reg_partial_sum(reg_psum_22_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_50( .activation_in(reg_activation_22_49), .weight_in(reg_weight_21_50), .partial_sum_in(reg_psum_21_50), .reg_activation(reg_activation_22_50), .reg_weight(reg_weight_22_50), .reg_partial_sum(reg_psum_22_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_51( .activation_in(reg_activation_22_50), .weight_in(reg_weight_21_51), .partial_sum_in(reg_psum_21_51), .reg_activation(reg_activation_22_51), .reg_weight(reg_weight_22_51), .reg_partial_sum(reg_psum_22_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_52( .activation_in(reg_activation_22_51), .weight_in(reg_weight_21_52), .partial_sum_in(reg_psum_21_52), .reg_activation(reg_activation_22_52), .reg_weight(reg_weight_22_52), .reg_partial_sum(reg_psum_22_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_53( .activation_in(reg_activation_22_52), .weight_in(reg_weight_21_53), .partial_sum_in(reg_psum_21_53), .reg_activation(reg_activation_22_53), .reg_weight(reg_weight_22_53), .reg_partial_sum(reg_psum_22_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_54( .activation_in(reg_activation_22_53), .weight_in(reg_weight_21_54), .partial_sum_in(reg_psum_21_54), .reg_activation(reg_activation_22_54), .reg_weight(reg_weight_22_54), .reg_partial_sum(reg_psum_22_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_55( .activation_in(reg_activation_22_54), .weight_in(reg_weight_21_55), .partial_sum_in(reg_psum_21_55), .reg_activation(reg_activation_22_55), .reg_weight(reg_weight_22_55), .reg_partial_sum(reg_psum_22_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_56( .activation_in(reg_activation_22_55), .weight_in(reg_weight_21_56), .partial_sum_in(reg_psum_21_56), .reg_activation(reg_activation_22_56), .reg_weight(reg_weight_22_56), .reg_partial_sum(reg_psum_22_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_57( .activation_in(reg_activation_22_56), .weight_in(reg_weight_21_57), .partial_sum_in(reg_psum_21_57), .reg_activation(reg_activation_22_57), .reg_weight(reg_weight_22_57), .reg_partial_sum(reg_psum_22_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_58( .activation_in(reg_activation_22_57), .weight_in(reg_weight_21_58), .partial_sum_in(reg_psum_21_58), .reg_activation(reg_activation_22_58), .reg_weight(reg_weight_22_58), .reg_partial_sum(reg_psum_22_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_59( .activation_in(reg_activation_22_58), .weight_in(reg_weight_21_59), .partial_sum_in(reg_psum_21_59), .reg_activation(reg_activation_22_59), .reg_weight(reg_weight_22_59), .reg_partial_sum(reg_psum_22_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_60( .activation_in(reg_activation_22_59), .weight_in(reg_weight_21_60), .partial_sum_in(reg_psum_21_60), .reg_activation(reg_activation_22_60), .reg_weight(reg_weight_22_60), .reg_partial_sum(reg_psum_22_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_61( .activation_in(reg_activation_22_60), .weight_in(reg_weight_21_61), .partial_sum_in(reg_psum_21_61), .reg_activation(reg_activation_22_61), .reg_weight(reg_weight_22_61), .reg_partial_sum(reg_psum_22_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_62( .activation_in(reg_activation_22_61), .weight_in(reg_weight_21_62), .partial_sum_in(reg_psum_21_62), .reg_activation(reg_activation_22_62), .reg_weight(reg_weight_22_62), .reg_partial_sum(reg_psum_22_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_63( .activation_in(reg_activation_22_62), .weight_in(reg_weight_21_63), .partial_sum_in(reg_psum_21_63), .reg_weight(reg_weight_22_63), .reg_partial_sum(reg_psum_22_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_0( .activation_in(in_activation_23), .weight_in(reg_weight_22_0), .partial_sum_in(reg_psum_22_0), .reg_activation(reg_activation_23_0), .reg_weight(reg_weight_23_0), .reg_partial_sum(reg_psum_23_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_1( .activation_in(reg_activation_23_0), .weight_in(reg_weight_22_1), .partial_sum_in(reg_psum_22_1), .reg_activation(reg_activation_23_1), .reg_weight(reg_weight_23_1), .reg_partial_sum(reg_psum_23_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_2( .activation_in(reg_activation_23_1), .weight_in(reg_weight_22_2), .partial_sum_in(reg_psum_22_2), .reg_activation(reg_activation_23_2), .reg_weight(reg_weight_23_2), .reg_partial_sum(reg_psum_23_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_3( .activation_in(reg_activation_23_2), .weight_in(reg_weight_22_3), .partial_sum_in(reg_psum_22_3), .reg_activation(reg_activation_23_3), .reg_weight(reg_weight_23_3), .reg_partial_sum(reg_psum_23_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_4( .activation_in(reg_activation_23_3), .weight_in(reg_weight_22_4), .partial_sum_in(reg_psum_22_4), .reg_activation(reg_activation_23_4), .reg_weight(reg_weight_23_4), .reg_partial_sum(reg_psum_23_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_5( .activation_in(reg_activation_23_4), .weight_in(reg_weight_22_5), .partial_sum_in(reg_psum_22_5), .reg_activation(reg_activation_23_5), .reg_weight(reg_weight_23_5), .reg_partial_sum(reg_psum_23_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_6( .activation_in(reg_activation_23_5), .weight_in(reg_weight_22_6), .partial_sum_in(reg_psum_22_6), .reg_activation(reg_activation_23_6), .reg_weight(reg_weight_23_6), .reg_partial_sum(reg_psum_23_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_7( .activation_in(reg_activation_23_6), .weight_in(reg_weight_22_7), .partial_sum_in(reg_psum_22_7), .reg_activation(reg_activation_23_7), .reg_weight(reg_weight_23_7), .reg_partial_sum(reg_psum_23_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_8( .activation_in(reg_activation_23_7), .weight_in(reg_weight_22_8), .partial_sum_in(reg_psum_22_8), .reg_activation(reg_activation_23_8), .reg_weight(reg_weight_23_8), .reg_partial_sum(reg_psum_23_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_9( .activation_in(reg_activation_23_8), .weight_in(reg_weight_22_9), .partial_sum_in(reg_psum_22_9), .reg_activation(reg_activation_23_9), .reg_weight(reg_weight_23_9), .reg_partial_sum(reg_psum_23_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_10( .activation_in(reg_activation_23_9), .weight_in(reg_weight_22_10), .partial_sum_in(reg_psum_22_10), .reg_activation(reg_activation_23_10), .reg_weight(reg_weight_23_10), .reg_partial_sum(reg_psum_23_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_11( .activation_in(reg_activation_23_10), .weight_in(reg_weight_22_11), .partial_sum_in(reg_psum_22_11), .reg_activation(reg_activation_23_11), .reg_weight(reg_weight_23_11), .reg_partial_sum(reg_psum_23_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_12( .activation_in(reg_activation_23_11), .weight_in(reg_weight_22_12), .partial_sum_in(reg_psum_22_12), .reg_activation(reg_activation_23_12), .reg_weight(reg_weight_23_12), .reg_partial_sum(reg_psum_23_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_13( .activation_in(reg_activation_23_12), .weight_in(reg_weight_22_13), .partial_sum_in(reg_psum_22_13), .reg_activation(reg_activation_23_13), .reg_weight(reg_weight_23_13), .reg_partial_sum(reg_psum_23_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_14( .activation_in(reg_activation_23_13), .weight_in(reg_weight_22_14), .partial_sum_in(reg_psum_22_14), .reg_activation(reg_activation_23_14), .reg_weight(reg_weight_23_14), .reg_partial_sum(reg_psum_23_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_15( .activation_in(reg_activation_23_14), .weight_in(reg_weight_22_15), .partial_sum_in(reg_psum_22_15), .reg_activation(reg_activation_23_15), .reg_weight(reg_weight_23_15), .reg_partial_sum(reg_psum_23_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_16( .activation_in(reg_activation_23_15), .weight_in(reg_weight_22_16), .partial_sum_in(reg_psum_22_16), .reg_activation(reg_activation_23_16), .reg_weight(reg_weight_23_16), .reg_partial_sum(reg_psum_23_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_17( .activation_in(reg_activation_23_16), .weight_in(reg_weight_22_17), .partial_sum_in(reg_psum_22_17), .reg_activation(reg_activation_23_17), .reg_weight(reg_weight_23_17), .reg_partial_sum(reg_psum_23_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_18( .activation_in(reg_activation_23_17), .weight_in(reg_weight_22_18), .partial_sum_in(reg_psum_22_18), .reg_activation(reg_activation_23_18), .reg_weight(reg_weight_23_18), .reg_partial_sum(reg_psum_23_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_19( .activation_in(reg_activation_23_18), .weight_in(reg_weight_22_19), .partial_sum_in(reg_psum_22_19), .reg_activation(reg_activation_23_19), .reg_weight(reg_weight_23_19), .reg_partial_sum(reg_psum_23_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_20( .activation_in(reg_activation_23_19), .weight_in(reg_weight_22_20), .partial_sum_in(reg_psum_22_20), .reg_activation(reg_activation_23_20), .reg_weight(reg_weight_23_20), .reg_partial_sum(reg_psum_23_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_21( .activation_in(reg_activation_23_20), .weight_in(reg_weight_22_21), .partial_sum_in(reg_psum_22_21), .reg_activation(reg_activation_23_21), .reg_weight(reg_weight_23_21), .reg_partial_sum(reg_psum_23_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_22( .activation_in(reg_activation_23_21), .weight_in(reg_weight_22_22), .partial_sum_in(reg_psum_22_22), .reg_activation(reg_activation_23_22), .reg_weight(reg_weight_23_22), .reg_partial_sum(reg_psum_23_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_23( .activation_in(reg_activation_23_22), .weight_in(reg_weight_22_23), .partial_sum_in(reg_psum_22_23), .reg_activation(reg_activation_23_23), .reg_weight(reg_weight_23_23), .reg_partial_sum(reg_psum_23_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_24( .activation_in(reg_activation_23_23), .weight_in(reg_weight_22_24), .partial_sum_in(reg_psum_22_24), .reg_activation(reg_activation_23_24), .reg_weight(reg_weight_23_24), .reg_partial_sum(reg_psum_23_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_25( .activation_in(reg_activation_23_24), .weight_in(reg_weight_22_25), .partial_sum_in(reg_psum_22_25), .reg_activation(reg_activation_23_25), .reg_weight(reg_weight_23_25), .reg_partial_sum(reg_psum_23_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_26( .activation_in(reg_activation_23_25), .weight_in(reg_weight_22_26), .partial_sum_in(reg_psum_22_26), .reg_activation(reg_activation_23_26), .reg_weight(reg_weight_23_26), .reg_partial_sum(reg_psum_23_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_27( .activation_in(reg_activation_23_26), .weight_in(reg_weight_22_27), .partial_sum_in(reg_psum_22_27), .reg_activation(reg_activation_23_27), .reg_weight(reg_weight_23_27), .reg_partial_sum(reg_psum_23_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_28( .activation_in(reg_activation_23_27), .weight_in(reg_weight_22_28), .partial_sum_in(reg_psum_22_28), .reg_activation(reg_activation_23_28), .reg_weight(reg_weight_23_28), .reg_partial_sum(reg_psum_23_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_29( .activation_in(reg_activation_23_28), .weight_in(reg_weight_22_29), .partial_sum_in(reg_psum_22_29), .reg_activation(reg_activation_23_29), .reg_weight(reg_weight_23_29), .reg_partial_sum(reg_psum_23_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_30( .activation_in(reg_activation_23_29), .weight_in(reg_weight_22_30), .partial_sum_in(reg_psum_22_30), .reg_activation(reg_activation_23_30), .reg_weight(reg_weight_23_30), .reg_partial_sum(reg_psum_23_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_31( .activation_in(reg_activation_23_30), .weight_in(reg_weight_22_31), .partial_sum_in(reg_psum_22_31), .reg_activation(reg_activation_23_31), .reg_weight(reg_weight_23_31), .reg_partial_sum(reg_psum_23_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_32( .activation_in(reg_activation_23_31), .weight_in(reg_weight_22_32), .partial_sum_in(reg_psum_22_32), .reg_activation(reg_activation_23_32), .reg_weight(reg_weight_23_32), .reg_partial_sum(reg_psum_23_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_33( .activation_in(reg_activation_23_32), .weight_in(reg_weight_22_33), .partial_sum_in(reg_psum_22_33), .reg_activation(reg_activation_23_33), .reg_weight(reg_weight_23_33), .reg_partial_sum(reg_psum_23_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_34( .activation_in(reg_activation_23_33), .weight_in(reg_weight_22_34), .partial_sum_in(reg_psum_22_34), .reg_activation(reg_activation_23_34), .reg_weight(reg_weight_23_34), .reg_partial_sum(reg_psum_23_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_35( .activation_in(reg_activation_23_34), .weight_in(reg_weight_22_35), .partial_sum_in(reg_psum_22_35), .reg_activation(reg_activation_23_35), .reg_weight(reg_weight_23_35), .reg_partial_sum(reg_psum_23_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_36( .activation_in(reg_activation_23_35), .weight_in(reg_weight_22_36), .partial_sum_in(reg_psum_22_36), .reg_activation(reg_activation_23_36), .reg_weight(reg_weight_23_36), .reg_partial_sum(reg_psum_23_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_37( .activation_in(reg_activation_23_36), .weight_in(reg_weight_22_37), .partial_sum_in(reg_psum_22_37), .reg_activation(reg_activation_23_37), .reg_weight(reg_weight_23_37), .reg_partial_sum(reg_psum_23_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_38( .activation_in(reg_activation_23_37), .weight_in(reg_weight_22_38), .partial_sum_in(reg_psum_22_38), .reg_activation(reg_activation_23_38), .reg_weight(reg_weight_23_38), .reg_partial_sum(reg_psum_23_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_39( .activation_in(reg_activation_23_38), .weight_in(reg_weight_22_39), .partial_sum_in(reg_psum_22_39), .reg_activation(reg_activation_23_39), .reg_weight(reg_weight_23_39), .reg_partial_sum(reg_psum_23_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_40( .activation_in(reg_activation_23_39), .weight_in(reg_weight_22_40), .partial_sum_in(reg_psum_22_40), .reg_activation(reg_activation_23_40), .reg_weight(reg_weight_23_40), .reg_partial_sum(reg_psum_23_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_41( .activation_in(reg_activation_23_40), .weight_in(reg_weight_22_41), .partial_sum_in(reg_psum_22_41), .reg_activation(reg_activation_23_41), .reg_weight(reg_weight_23_41), .reg_partial_sum(reg_psum_23_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_42( .activation_in(reg_activation_23_41), .weight_in(reg_weight_22_42), .partial_sum_in(reg_psum_22_42), .reg_activation(reg_activation_23_42), .reg_weight(reg_weight_23_42), .reg_partial_sum(reg_psum_23_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_43( .activation_in(reg_activation_23_42), .weight_in(reg_weight_22_43), .partial_sum_in(reg_psum_22_43), .reg_activation(reg_activation_23_43), .reg_weight(reg_weight_23_43), .reg_partial_sum(reg_psum_23_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_44( .activation_in(reg_activation_23_43), .weight_in(reg_weight_22_44), .partial_sum_in(reg_psum_22_44), .reg_activation(reg_activation_23_44), .reg_weight(reg_weight_23_44), .reg_partial_sum(reg_psum_23_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_45( .activation_in(reg_activation_23_44), .weight_in(reg_weight_22_45), .partial_sum_in(reg_psum_22_45), .reg_activation(reg_activation_23_45), .reg_weight(reg_weight_23_45), .reg_partial_sum(reg_psum_23_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_46( .activation_in(reg_activation_23_45), .weight_in(reg_weight_22_46), .partial_sum_in(reg_psum_22_46), .reg_activation(reg_activation_23_46), .reg_weight(reg_weight_23_46), .reg_partial_sum(reg_psum_23_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_47( .activation_in(reg_activation_23_46), .weight_in(reg_weight_22_47), .partial_sum_in(reg_psum_22_47), .reg_activation(reg_activation_23_47), .reg_weight(reg_weight_23_47), .reg_partial_sum(reg_psum_23_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_48( .activation_in(reg_activation_23_47), .weight_in(reg_weight_22_48), .partial_sum_in(reg_psum_22_48), .reg_activation(reg_activation_23_48), .reg_weight(reg_weight_23_48), .reg_partial_sum(reg_psum_23_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_49( .activation_in(reg_activation_23_48), .weight_in(reg_weight_22_49), .partial_sum_in(reg_psum_22_49), .reg_activation(reg_activation_23_49), .reg_weight(reg_weight_23_49), .reg_partial_sum(reg_psum_23_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_50( .activation_in(reg_activation_23_49), .weight_in(reg_weight_22_50), .partial_sum_in(reg_psum_22_50), .reg_activation(reg_activation_23_50), .reg_weight(reg_weight_23_50), .reg_partial_sum(reg_psum_23_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_51( .activation_in(reg_activation_23_50), .weight_in(reg_weight_22_51), .partial_sum_in(reg_psum_22_51), .reg_activation(reg_activation_23_51), .reg_weight(reg_weight_23_51), .reg_partial_sum(reg_psum_23_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_52( .activation_in(reg_activation_23_51), .weight_in(reg_weight_22_52), .partial_sum_in(reg_psum_22_52), .reg_activation(reg_activation_23_52), .reg_weight(reg_weight_23_52), .reg_partial_sum(reg_psum_23_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_53( .activation_in(reg_activation_23_52), .weight_in(reg_weight_22_53), .partial_sum_in(reg_psum_22_53), .reg_activation(reg_activation_23_53), .reg_weight(reg_weight_23_53), .reg_partial_sum(reg_psum_23_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_54( .activation_in(reg_activation_23_53), .weight_in(reg_weight_22_54), .partial_sum_in(reg_psum_22_54), .reg_activation(reg_activation_23_54), .reg_weight(reg_weight_23_54), .reg_partial_sum(reg_psum_23_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_55( .activation_in(reg_activation_23_54), .weight_in(reg_weight_22_55), .partial_sum_in(reg_psum_22_55), .reg_activation(reg_activation_23_55), .reg_weight(reg_weight_23_55), .reg_partial_sum(reg_psum_23_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_56( .activation_in(reg_activation_23_55), .weight_in(reg_weight_22_56), .partial_sum_in(reg_psum_22_56), .reg_activation(reg_activation_23_56), .reg_weight(reg_weight_23_56), .reg_partial_sum(reg_psum_23_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_57( .activation_in(reg_activation_23_56), .weight_in(reg_weight_22_57), .partial_sum_in(reg_psum_22_57), .reg_activation(reg_activation_23_57), .reg_weight(reg_weight_23_57), .reg_partial_sum(reg_psum_23_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_58( .activation_in(reg_activation_23_57), .weight_in(reg_weight_22_58), .partial_sum_in(reg_psum_22_58), .reg_activation(reg_activation_23_58), .reg_weight(reg_weight_23_58), .reg_partial_sum(reg_psum_23_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_59( .activation_in(reg_activation_23_58), .weight_in(reg_weight_22_59), .partial_sum_in(reg_psum_22_59), .reg_activation(reg_activation_23_59), .reg_weight(reg_weight_23_59), .reg_partial_sum(reg_psum_23_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_60( .activation_in(reg_activation_23_59), .weight_in(reg_weight_22_60), .partial_sum_in(reg_psum_22_60), .reg_activation(reg_activation_23_60), .reg_weight(reg_weight_23_60), .reg_partial_sum(reg_psum_23_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_61( .activation_in(reg_activation_23_60), .weight_in(reg_weight_22_61), .partial_sum_in(reg_psum_22_61), .reg_activation(reg_activation_23_61), .reg_weight(reg_weight_23_61), .reg_partial_sum(reg_psum_23_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_62( .activation_in(reg_activation_23_61), .weight_in(reg_weight_22_62), .partial_sum_in(reg_psum_22_62), .reg_activation(reg_activation_23_62), .reg_weight(reg_weight_23_62), .reg_partial_sum(reg_psum_23_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_63( .activation_in(reg_activation_23_62), .weight_in(reg_weight_22_63), .partial_sum_in(reg_psum_22_63), .reg_weight(reg_weight_23_63), .reg_partial_sum(reg_psum_23_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_0( .activation_in(in_activation_24), .weight_in(reg_weight_23_0), .partial_sum_in(reg_psum_23_0), .reg_activation(reg_activation_24_0), .reg_weight(reg_weight_24_0), .reg_partial_sum(reg_psum_24_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_1( .activation_in(reg_activation_24_0), .weight_in(reg_weight_23_1), .partial_sum_in(reg_psum_23_1), .reg_activation(reg_activation_24_1), .reg_weight(reg_weight_24_1), .reg_partial_sum(reg_psum_24_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_2( .activation_in(reg_activation_24_1), .weight_in(reg_weight_23_2), .partial_sum_in(reg_psum_23_2), .reg_activation(reg_activation_24_2), .reg_weight(reg_weight_24_2), .reg_partial_sum(reg_psum_24_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_3( .activation_in(reg_activation_24_2), .weight_in(reg_weight_23_3), .partial_sum_in(reg_psum_23_3), .reg_activation(reg_activation_24_3), .reg_weight(reg_weight_24_3), .reg_partial_sum(reg_psum_24_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_4( .activation_in(reg_activation_24_3), .weight_in(reg_weight_23_4), .partial_sum_in(reg_psum_23_4), .reg_activation(reg_activation_24_4), .reg_weight(reg_weight_24_4), .reg_partial_sum(reg_psum_24_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_5( .activation_in(reg_activation_24_4), .weight_in(reg_weight_23_5), .partial_sum_in(reg_psum_23_5), .reg_activation(reg_activation_24_5), .reg_weight(reg_weight_24_5), .reg_partial_sum(reg_psum_24_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_6( .activation_in(reg_activation_24_5), .weight_in(reg_weight_23_6), .partial_sum_in(reg_psum_23_6), .reg_activation(reg_activation_24_6), .reg_weight(reg_weight_24_6), .reg_partial_sum(reg_psum_24_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_7( .activation_in(reg_activation_24_6), .weight_in(reg_weight_23_7), .partial_sum_in(reg_psum_23_7), .reg_activation(reg_activation_24_7), .reg_weight(reg_weight_24_7), .reg_partial_sum(reg_psum_24_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_8( .activation_in(reg_activation_24_7), .weight_in(reg_weight_23_8), .partial_sum_in(reg_psum_23_8), .reg_activation(reg_activation_24_8), .reg_weight(reg_weight_24_8), .reg_partial_sum(reg_psum_24_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_9( .activation_in(reg_activation_24_8), .weight_in(reg_weight_23_9), .partial_sum_in(reg_psum_23_9), .reg_activation(reg_activation_24_9), .reg_weight(reg_weight_24_9), .reg_partial_sum(reg_psum_24_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_10( .activation_in(reg_activation_24_9), .weight_in(reg_weight_23_10), .partial_sum_in(reg_psum_23_10), .reg_activation(reg_activation_24_10), .reg_weight(reg_weight_24_10), .reg_partial_sum(reg_psum_24_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_11( .activation_in(reg_activation_24_10), .weight_in(reg_weight_23_11), .partial_sum_in(reg_psum_23_11), .reg_activation(reg_activation_24_11), .reg_weight(reg_weight_24_11), .reg_partial_sum(reg_psum_24_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_12( .activation_in(reg_activation_24_11), .weight_in(reg_weight_23_12), .partial_sum_in(reg_psum_23_12), .reg_activation(reg_activation_24_12), .reg_weight(reg_weight_24_12), .reg_partial_sum(reg_psum_24_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_13( .activation_in(reg_activation_24_12), .weight_in(reg_weight_23_13), .partial_sum_in(reg_psum_23_13), .reg_activation(reg_activation_24_13), .reg_weight(reg_weight_24_13), .reg_partial_sum(reg_psum_24_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_14( .activation_in(reg_activation_24_13), .weight_in(reg_weight_23_14), .partial_sum_in(reg_psum_23_14), .reg_activation(reg_activation_24_14), .reg_weight(reg_weight_24_14), .reg_partial_sum(reg_psum_24_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_15( .activation_in(reg_activation_24_14), .weight_in(reg_weight_23_15), .partial_sum_in(reg_psum_23_15), .reg_activation(reg_activation_24_15), .reg_weight(reg_weight_24_15), .reg_partial_sum(reg_psum_24_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_16( .activation_in(reg_activation_24_15), .weight_in(reg_weight_23_16), .partial_sum_in(reg_psum_23_16), .reg_activation(reg_activation_24_16), .reg_weight(reg_weight_24_16), .reg_partial_sum(reg_psum_24_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_17( .activation_in(reg_activation_24_16), .weight_in(reg_weight_23_17), .partial_sum_in(reg_psum_23_17), .reg_activation(reg_activation_24_17), .reg_weight(reg_weight_24_17), .reg_partial_sum(reg_psum_24_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_18( .activation_in(reg_activation_24_17), .weight_in(reg_weight_23_18), .partial_sum_in(reg_psum_23_18), .reg_activation(reg_activation_24_18), .reg_weight(reg_weight_24_18), .reg_partial_sum(reg_psum_24_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_19( .activation_in(reg_activation_24_18), .weight_in(reg_weight_23_19), .partial_sum_in(reg_psum_23_19), .reg_activation(reg_activation_24_19), .reg_weight(reg_weight_24_19), .reg_partial_sum(reg_psum_24_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_20( .activation_in(reg_activation_24_19), .weight_in(reg_weight_23_20), .partial_sum_in(reg_psum_23_20), .reg_activation(reg_activation_24_20), .reg_weight(reg_weight_24_20), .reg_partial_sum(reg_psum_24_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_21( .activation_in(reg_activation_24_20), .weight_in(reg_weight_23_21), .partial_sum_in(reg_psum_23_21), .reg_activation(reg_activation_24_21), .reg_weight(reg_weight_24_21), .reg_partial_sum(reg_psum_24_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_22( .activation_in(reg_activation_24_21), .weight_in(reg_weight_23_22), .partial_sum_in(reg_psum_23_22), .reg_activation(reg_activation_24_22), .reg_weight(reg_weight_24_22), .reg_partial_sum(reg_psum_24_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_23( .activation_in(reg_activation_24_22), .weight_in(reg_weight_23_23), .partial_sum_in(reg_psum_23_23), .reg_activation(reg_activation_24_23), .reg_weight(reg_weight_24_23), .reg_partial_sum(reg_psum_24_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_24( .activation_in(reg_activation_24_23), .weight_in(reg_weight_23_24), .partial_sum_in(reg_psum_23_24), .reg_activation(reg_activation_24_24), .reg_weight(reg_weight_24_24), .reg_partial_sum(reg_psum_24_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_25( .activation_in(reg_activation_24_24), .weight_in(reg_weight_23_25), .partial_sum_in(reg_psum_23_25), .reg_activation(reg_activation_24_25), .reg_weight(reg_weight_24_25), .reg_partial_sum(reg_psum_24_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_26( .activation_in(reg_activation_24_25), .weight_in(reg_weight_23_26), .partial_sum_in(reg_psum_23_26), .reg_activation(reg_activation_24_26), .reg_weight(reg_weight_24_26), .reg_partial_sum(reg_psum_24_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_27( .activation_in(reg_activation_24_26), .weight_in(reg_weight_23_27), .partial_sum_in(reg_psum_23_27), .reg_activation(reg_activation_24_27), .reg_weight(reg_weight_24_27), .reg_partial_sum(reg_psum_24_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_28( .activation_in(reg_activation_24_27), .weight_in(reg_weight_23_28), .partial_sum_in(reg_psum_23_28), .reg_activation(reg_activation_24_28), .reg_weight(reg_weight_24_28), .reg_partial_sum(reg_psum_24_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_29( .activation_in(reg_activation_24_28), .weight_in(reg_weight_23_29), .partial_sum_in(reg_psum_23_29), .reg_activation(reg_activation_24_29), .reg_weight(reg_weight_24_29), .reg_partial_sum(reg_psum_24_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_30( .activation_in(reg_activation_24_29), .weight_in(reg_weight_23_30), .partial_sum_in(reg_psum_23_30), .reg_activation(reg_activation_24_30), .reg_weight(reg_weight_24_30), .reg_partial_sum(reg_psum_24_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_31( .activation_in(reg_activation_24_30), .weight_in(reg_weight_23_31), .partial_sum_in(reg_psum_23_31), .reg_activation(reg_activation_24_31), .reg_weight(reg_weight_24_31), .reg_partial_sum(reg_psum_24_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_32( .activation_in(reg_activation_24_31), .weight_in(reg_weight_23_32), .partial_sum_in(reg_psum_23_32), .reg_activation(reg_activation_24_32), .reg_weight(reg_weight_24_32), .reg_partial_sum(reg_psum_24_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_33( .activation_in(reg_activation_24_32), .weight_in(reg_weight_23_33), .partial_sum_in(reg_psum_23_33), .reg_activation(reg_activation_24_33), .reg_weight(reg_weight_24_33), .reg_partial_sum(reg_psum_24_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_34( .activation_in(reg_activation_24_33), .weight_in(reg_weight_23_34), .partial_sum_in(reg_psum_23_34), .reg_activation(reg_activation_24_34), .reg_weight(reg_weight_24_34), .reg_partial_sum(reg_psum_24_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_35( .activation_in(reg_activation_24_34), .weight_in(reg_weight_23_35), .partial_sum_in(reg_psum_23_35), .reg_activation(reg_activation_24_35), .reg_weight(reg_weight_24_35), .reg_partial_sum(reg_psum_24_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_36( .activation_in(reg_activation_24_35), .weight_in(reg_weight_23_36), .partial_sum_in(reg_psum_23_36), .reg_activation(reg_activation_24_36), .reg_weight(reg_weight_24_36), .reg_partial_sum(reg_psum_24_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_37( .activation_in(reg_activation_24_36), .weight_in(reg_weight_23_37), .partial_sum_in(reg_psum_23_37), .reg_activation(reg_activation_24_37), .reg_weight(reg_weight_24_37), .reg_partial_sum(reg_psum_24_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_38( .activation_in(reg_activation_24_37), .weight_in(reg_weight_23_38), .partial_sum_in(reg_psum_23_38), .reg_activation(reg_activation_24_38), .reg_weight(reg_weight_24_38), .reg_partial_sum(reg_psum_24_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_39( .activation_in(reg_activation_24_38), .weight_in(reg_weight_23_39), .partial_sum_in(reg_psum_23_39), .reg_activation(reg_activation_24_39), .reg_weight(reg_weight_24_39), .reg_partial_sum(reg_psum_24_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_40( .activation_in(reg_activation_24_39), .weight_in(reg_weight_23_40), .partial_sum_in(reg_psum_23_40), .reg_activation(reg_activation_24_40), .reg_weight(reg_weight_24_40), .reg_partial_sum(reg_psum_24_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_41( .activation_in(reg_activation_24_40), .weight_in(reg_weight_23_41), .partial_sum_in(reg_psum_23_41), .reg_activation(reg_activation_24_41), .reg_weight(reg_weight_24_41), .reg_partial_sum(reg_psum_24_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_42( .activation_in(reg_activation_24_41), .weight_in(reg_weight_23_42), .partial_sum_in(reg_psum_23_42), .reg_activation(reg_activation_24_42), .reg_weight(reg_weight_24_42), .reg_partial_sum(reg_psum_24_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_43( .activation_in(reg_activation_24_42), .weight_in(reg_weight_23_43), .partial_sum_in(reg_psum_23_43), .reg_activation(reg_activation_24_43), .reg_weight(reg_weight_24_43), .reg_partial_sum(reg_psum_24_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_44( .activation_in(reg_activation_24_43), .weight_in(reg_weight_23_44), .partial_sum_in(reg_psum_23_44), .reg_activation(reg_activation_24_44), .reg_weight(reg_weight_24_44), .reg_partial_sum(reg_psum_24_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_45( .activation_in(reg_activation_24_44), .weight_in(reg_weight_23_45), .partial_sum_in(reg_psum_23_45), .reg_activation(reg_activation_24_45), .reg_weight(reg_weight_24_45), .reg_partial_sum(reg_psum_24_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_46( .activation_in(reg_activation_24_45), .weight_in(reg_weight_23_46), .partial_sum_in(reg_psum_23_46), .reg_activation(reg_activation_24_46), .reg_weight(reg_weight_24_46), .reg_partial_sum(reg_psum_24_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_47( .activation_in(reg_activation_24_46), .weight_in(reg_weight_23_47), .partial_sum_in(reg_psum_23_47), .reg_activation(reg_activation_24_47), .reg_weight(reg_weight_24_47), .reg_partial_sum(reg_psum_24_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_48( .activation_in(reg_activation_24_47), .weight_in(reg_weight_23_48), .partial_sum_in(reg_psum_23_48), .reg_activation(reg_activation_24_48), .reg_weight(reg_weight_24_48), .reg_partial_sum(reg_psum_24_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_49( .activation_in(reg_activation_24_48), .weight_in(reg_weight_23_49), .partial_sum_in(reg_psum_23_49), .reg_activation(reg_activation_24_49), .reg_weight(reg_weight_24_49), .reg_partial_sum(reg_psum_24_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_50( .activation_in(reg_activation_24_49), .weight_in(reg_weight_23_50), .partial_sum_in(reg_psum_23_50), .reg_activation(reg_activation_24_50), .reg_weight(reg_weight_24_50), .reg_partial_sum(reg_psum_24_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_51( .activation_in(reg_activation_24_50), .weight_in(reg_weight_23_51), .partial_sum_in(reg_psum_23_51), .reg_activation(reg_activation_24_51), .reg_weight(reg_weight_24_51), .reg_partial_sum(reg_psum_24_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_52( .activation_in(reg_activation_24_51), .weight_in(reg_weight_23_52), .partial_sum_in(reg_psum_23_52), .reg_activation(reg_activation_24_52), .reg_weight(reg_weight_24_52), .reg_partial_sum(reg_psum_24_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_53( .activation_in(reg_activation_24_52), .weight_in(reg_weight_23_53), .partial_sum_in(reg_psum_23_53), .reg_activation(reg_activation_24_53), .reg_weight(reg_weight_24_53), .reg_partial_sum(reg_psum_24_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_54( .activation_in(reg_activation_24_53), .weight_in(reg_weight_23_54), .partial_sum_in(reg_psum_23_54), .reg_activation(reg_activation_24_54), .reg_weight(reg_weight_24_54), .reg_partial_sum(reg_psum_24_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_55( .activation_in(reg_activation_24_54), .weight_in(reg_weight_23_55), .partial_sum_in(reg_psum_23_55), .reg_activation(reg_activation_24_55), .reg_weight(reg_weight_24_55), .reg_partial_sum(reg_psum_24_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_56( .activation_in(reg_activation_24_55), .weight_in(reg_weight_23_56), .partial_sum_in(reg_psum_23_56), .reg_activation(reg_activation_24_56), .reg_weight(reg_weight_24_56), .reg_partial_sum(reg_psum_24_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_57( .activation_in(reg_activation_24_56), .weight_in(reg_weight_23_57), .partial_sum_in(reg_psum_23_57), .reg_activation(reg_activation_24_57), .reg_weight(reg_weight_24_57), .reg_partial_sum(reg_psum_24_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_58( .activation_in(reg_activation_24_57), .weight_in(reg_weight_23_58), .partial_sum_in(reg_psum_23_58), .reg_activation(reg_activation_24_58), .reg_weight(reg_weight_24_58), .reg_partial_sum(reg_psum_24_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_59( .activation_in(reg_activation_24_58), .weight_in(reg_weight_23_59), .partial_sum_in(reg_psum_23_59), .reg_activation(reg_activation_24_59), .reg_weight(reg_weight_24_59), .reg_partial_sum(reg_psum_24_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_60( .activation_in(reg_activation_24_59), .weight_in(reg_weight_23_60), .partial_sum_in(reg_psum_23_60), .reg_activation(reg_activation_24_60), .reg_weight(reg_weight_24_60), .reg_partial_sum(reg_psum_24_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_61( .activation_in(reg_activation_24_60), .weight_in(reg_weight_23_61), .partial_sum_in(reg_psum_23_61), .reg_activation(reg_activation_24_61), .reg_weight(reg_weight_24_61), .reg_partial_sum(reg_psum_24_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_62( .activation_in(reg_activation_24_61), .weight_in(reg_weight_23_62), .partial_sum_in(reg_psum_23_62), .reg_activation(reg_activation_24_62), .reg_weight(reg_weight_24_62), .reg_partial_sum(reg_psum_24_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_63( .activation_in(reg_activation_24_62), .weight_in(reg_weight_23_63), .partial_sum_in(reg_psum_23_63), .reg_weight(reg_weight_24_63), .reg_partial_sum(reg_psum_24_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_0( .activation_in(in_activation_25), .weight_in(reg_weight_24_0), .partial_sum_in(reg_psum_24_0), .reg_activation(reg_activation_25_0), .reg_weight(reg_weight_25_0), .reg_partial_sum(reg_psum_25_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_1( .activation_in(reg_activation_25_0), .weight_in(reg_weight_24_1), .partial_sum_in(reg_psum_24_1), .reg_activation(reg_activation_25_1), .reg_weight(reg_weight_25_1), .reg_partial_sum(reg_psum_25_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_2( .activation_in(reg_activation_25_1), .weight_in(reg_weight_24_2), .partial_sum_in(reg_psum_24_2), .reg_activation(reg_activation_25_2), .reg_weight(reg_weight_25_2), .reg_partial_sum(reg_psum_25_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_3( .activation_in(reg_activation_25_2), .weight_in(reg_weight_24_3), .partial_sum_in(reg_psum_24_3), .reg_activation(reg_activation_25_3), .reg_weight(reg_weight_25_3), .reg_partial_sum(reg_psum_25_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_4( .activation_in(reg_activation_25_3), .weight_in(reg_weight_24_4), .partial_sum_in(reg_psum_24_4), .reg_activation(reg_activation_25_4), .reg_weight(reg_weight_25_4), .reg_partial_sum(reg_psum_25_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_5( .activation_in(reg_activation_25_4), .weight_in(reg_weight_24_5), .partial_sum_in(reg_psum_24_5), .reg_activation(reg_activation_25_5), .reg_weight(reg_weight_25_5), .reg_partial_sum(reg_psum_25_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_6( .activation_in(reg_activation_25_5), .weight_in(reg_weight_24_6), .partial_sum_in(reg_psum_24_6), .reg_activation(reg_activation_25_6), .reg_weight(reg_weight_25_6), .reg_partial_sum(reg_psum_25_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_7( .activation_in(reg_activation_25_6), .weight_in(reg_weight_24_7), .partial_sum_in(reg_psum_24_7), .reg_activation(reg_activation_25_7), .reg_weight(reg_weight_25_7), .reg_partial_sum(reg_psum_25_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_8( .activation_in(reg_activation_25_7), .weight_in(reg_weight_24_8), .partial_sum_in(reg_psum_24_8), .reg_activation(reg_activation_25_8), .reg_weight(reg_weight_25_8), .reg_partial_sum(reg_psum_25_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_9( .activation_in(reg_activation_25_8), .weight_in(reg_weight_24_9), .partial_sum_in(reg_psum_24_9), .reg_activation(reg_activation_25_9), .reg_weight(reg_weight_25_9), .reg_partial_sum(reg_psum_25_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_10( .activation_in(reg_activation_25_9), .weight_in(reg_weight_24_10), .partial_sum_in(reg_psum_24_10), .reg_activation(reg_activation_25_10), .reg_weight(reg_weight_25_10), .reg_partial_sum(reg_psum_25_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_11( .activation_in(reg_activation_25_10), .weight_in(reg_weight_24_11), .partial_sum_in(reg_psum_24_11), .reg_activation(reg_activation_25_11), .reg_weight(reg_weight_25_11), .reg_partial_sum(reg_psum_25_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_12( .activation_in(reg_activation_25_11), .weight_in(reg_weight_24_12), .partial_sum_in(reg_psum_24_12), .reg_activation(reg_activation_25_12), .reg_weight(reg_weight_25_12), .reg_partial_sum(reg_psum_25_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_13( .activation_in(reg_activation_25_12), .weight_in(reg_weight_24_13), .partial_sum_in(reg_psum_24_13), .reg_activation(reg_activation_25_13), .reg_weight(reg_weight_25_13), .reg_partial_sum(reg_psum_25_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_14( .activation_in(reg_activation_25_13), .weight_in(reg_weight_24_14), .partial_sum_in(reg_psum_24_14), .reg_activation(reg_activation_25_14), .reg_weight(reg_weight_25_14), .reg_partial_sum(reg_psum_25_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_15( .activation_in(reg_activation_25_14), .weight_in(reg_weight_24_15), .partial_sum_in(reg_psum_24_15), .reg_activation(reg_activation_25_15), .reg_weight(reg_weight_25_15), .reg_partial_sum(reg_psum_25_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_16( .activation_in(reg_activation_25_15), .weight_in(reg_weight_24_16), .partial_sum_in(reg_psum_24_16), .reg_activation(reg_activation_25_16), .reg_weight(reg_weight_25_16), .reg_partial_sum(reg_psum_25_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_17( .activation_in(reg_activation_25_16), .weight_in(reg_weight_24_17), .partial_sum_in(reg_psum_24_17), .reg_activation(reg_activation_25_17), .reg_weight(reg_weight_25_17), .reg_partial_sum(reg_psum_25_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_18( .activation_in(reg_activation_25_17), .weight_in(reg_weight_24_18), .partial_sum_in(reg_psum_24_18), .reg_activation(reg_activation_25_18), .reg_weight(reg_weight_25_18), .reg_partial_sum(reg_psum_25_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_19( .activation_in(reg_activation_25_18), .weight_in(reg_weight_24_19), .partial_sum_in(reg_psum_24_19), .reg_activation(reg_activation_25_19), .reg_weight(reg_weight_25_19), .reg_partial_sum(reg_psum_25_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_20( .activation_in(reg_activation_25_19), .weight_in(reg_weight_24_20), .partial_sum_in(reg_psum_24_20), .reg_activation(reg_activation_25_20), .reg_weight(reg_weight_25_20), .reg_partial_sum(reg_psum_25_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_21( .activation_in(reg_activation_25_20), .weight_in(reg_weight_24_21), .partial_sum_in(reg_psum_24_21), .reg_activation(reg_activation_25_21), .reg_weight(reg_weight_25_21), .reg_partial_sum(reg_psum_25_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_22( .activation_in(reg_activation_25_21), .weight_in(reg_weight_24_22), .partial_sum_in(reg_psum_24_22), .reg_activation(reg_activation_25_22), .reg_weight(reg_weight_25_22), .reg_partial_sum(reg_psum_25_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_23( .activation_in(reg_activation_25_22), .weight_in(reg_weight_24_23), .partial_sum_in(reg_psum_24_23), .reg_activation(reg_activation_25_23), .reg_weight(reg_weight_25_23), .reg_partial_sum(reg_psum_25_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_24( .activation_in(reg_activation_25_23), .weight_in(reg_weight_24_24), .partial_sum_in(reg_psum_24_24), .reg_activation(reg_activation_25_24), .reg_weight(reg_weight_25_24), .reg_partial_sum(reg_psum_25_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_25( .activation_in(reg_activation_25_24), .weight_in(reg_weight_24_25), .partial_sum_in(reg_psum_24_25), .reg_activation(reg_activation_25_25), .reg_weight(reg_weight_25_25), .reg_partial_sum(reg_psum_25_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_26( .activation_in(reg_activation_25_25), .weight_in(reg_weight_24_26), .partial_sum_in(reg_psum_24_26), .reg_activation(reg_activation_25_26), .reg_weight(reg_weight_25_26), .reg_partial_sum(reg_psum_25_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_27( .activation_in(reg_activation_25_26), .weight_in(reg_weight_24_27), .partial_sum_in(reg_psum_24_27), .reg_activation(reg_activation_25_27), .reg_weight(reg_weight_25_27), .reg_partial_sum(reg_psum_25_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_28( .activation_in(reg_activation_25_27), .weight_in(reg_weight_24_28), .partial_sum_in(reg_psum_24_28), .reg_activation(reg_activation_25_28), .reg_weight(reg_weight_25_28), .reg_partial_sum(reg_psum_25_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_29( .activation_in(reg_activation_25_28), .weight_in(reg_weight_24_29), .partial_sum_in(reg_psum_24_29), .reg_activation(reg_activation_25_29), .reg_weight(reg_weight_25_29), .reg_partial_sum(reg_psum_25_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_30( .activation_in(reg_activation_25_29), .weight_in(reg_weight_24_30), .partial_sum_in(reg_psum_24_30), .reg_activation(reg_activation_25_30), .reg_weight(reg_weight_25_30), .reg_partial_sum(reg_psum_25_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_31( .activation_in(reg_activation_25_30), .weight_in(reg_weight_24_31), .partial_sum_in(reg_psum_24_31), .reg_activation(reg_activation_25_31), .reg_weight(reg_weight_25_31), .reg_partial_sum(reg_psum_25_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_32( .activation_in(reg_activation_25_31), .weight_in(reg_weight_24_32), .partial_sum_in(reg_psum_24_32), .reg_activation(reg_activation_25_32), .reg_weight(reg_weight_25_32), .reg_partial_sum(reg_psum_25_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_33( .activation_in(reg_activation_25_32), .weight_in(reg_weight_24_33), .partial_sum_in(reg_psum_24_33), .reg_activation(reg_activation_25_33), .reg_weight(reg_weight_25_33), .reg_partial_sum(reg_psum_25_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_34( .activation_in(reg_activation_25_33), .weight_in(reg_weight_24_34), .partial_sum_in(reg_psum_24_34), .reg_activation(reg_activation_25_34), .reg_weight(reg_weight_25_34), .reg_partial_sum(reg_psum_25_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_35( .activation_in(reg_activation_25_34), .weight_in(reg_weight_24_35), .partial_sum_in(reg_psum_24_35), .reg_activation(reg_activation_25_35), .reg_weight(reg_weight_25_35), .reg_partial_sum(reg_psum_25_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_36( .activation_in(reg_activation_25_35), .weight_in(reg_weight_24_36), .partial_sum_in(reg_psum_24_36), .reg_activation(reg_activation_25_36), .reg_weight(reg_weight_25_36), .reg_partial_sum(reg_psum_25_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_37( .activation_in(reg_activation_25_36), .weight_in(reg_weight_24_37), .partial_sum_in(reg_psum_24_37), .reg_activation(reg_activation_25_37), .reg_weight(reg_weight_25_37), .reg_partial_sum(reg_psum_25_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_38( .activation_in(reg_activation_25_37), .weight_in(reg_weight_24_38), .partial_sum_in(reg_psum_24_38), .reg_activation(reg_activation_25_38), .reg_weight(reg_weight_25_38), .reg_partial_sum(reg_psum_25_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_39( .activation_in(reg_activation_25_38), .weight_in(reg_weight_24_39), .partial_sum_in(reg_psum_24_39), .reg_activation(reg_activation_25_39), .reg_weight(reg_weight_25_39), .reg_partial_sum(reg_psum_25_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_40( .activation_in(reg_activation_25_39), .weight_in(reg_weight_24_40), .partial_sum_in(reg_psum_24_40), .reg_activation(reg_activation_25_40), .reg_weight(reg_weight_25_40), .reg_partial_sum(reg_psum_25_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_41( .activation_in(reg_activation_25_40), .weight_in(reg_weight_24_41), .partial_sum_in(reg_psum_24_41), .reg_activation(reg_activation_25_41), .reg_weight(reg_weight_25_41), .reg_partial_sum(reg_psum_25_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_42( .activation_in(reg_activation_25_41), .weight_in(reg_weight_24_42), .partial_sum_in(reg_psum_24_42), .reg_activation(reg_activation_25_42), .reg_weight(reg_weight_25_42), .reg_partial_sum(reg_psum_25_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_43( .activation_in(reg_activation_25_42), .weight_in(reg_weight_24_43), .partial_sum_in(reg_psum_24_43), .reg_activation(reg_activation_25_43), .reg_weight(reg_weight_25_43), .reg_partial_sum(reg_psum_25_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_44( .activation_in(reg_activation_25_43), .weight_in(reg_weight_24_44), .partial_sum_in(reg_psum_24_44), .reg_activation(reg_activation_25_44), .reg_weight(reg_weight_25_44), .reg_partial_sum(reg_psum_25_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_45( .activation_in(reg_activation_25_44), .weight_in(reg_weight_24_45), .partial_sum_in(reg_psum_24_45), .reg_activation(reg_activation_25_45), .reg_weight(reg_weight_25_45), .reg_partial_sum(reg_psum_25_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_46( .activation_in(reg_activation_25_45), .weight_in(reg_weight_24_46), .partial_sum_in(reg_psum_24_46), .reg_activation(reg_activation_25_46), .reg_weight(reg_weight_25_46), .reg_partial_sum(reg_psum_25_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_47( .activation_in(reg_activation_25_46), .weight_in(reg_weight_24_47), .partial_sum_in(reg_psum_24_47), .reg_activation(reg_activation_25_47), .reg_weight(reg_weight_25_47), .reg_partial_sum(reg_psum_25_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_48( .activation_in(reg_activation_25_47), .weight_in(reg_weight_24_48), .partial_sum_in(reg_psum_24_48), .reg_activation(reg_activation_25_48), .reg_weight(reg_weight_25_48), .reg_partial_sum(reg_psum_25_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_49( .activation_in(reg_activation_25_48), .weight_in(reg_weight_24_49), .partial_sum_in(reg_psum_24_49), .reg_activation(reg_activation_25_49), .reg_weight(reg_weight_25_49), .reg_partial_sum(reg_psum_25_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_50( .activation_in(reg_activation_25_49), .weight_in(reg_weight_24_50), .partial_sum_in(reg_psum_24_50), .reg_activation(reg_activation_25_50), .reg_weight(reg_weight_25_50), .reg_partial_sum(reg_psum_25_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_51( .activation_in(reg_activation_25_50), .weight_in(reg_weight_24_51), .partial_sum_in(reg_psum_24_51), .reg_activation(reg_activation_25_51), .reg_weight(reg_weight_25_51), .reg_partial_sum(reg_psum_25_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_52( .activation_in(reg_activation_25_51), .weight_in(reg_weight_24_52), .partial_sum_in(reg_psum_24_52), .reg_activation(reg_activation_25_52), .reg_weight(reg_weight_25_52), .reg_partial_sum(reg_psum_25_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_53( .activation_in(reg_activation_25_52), .weight_in(reg_weight_24_53), .partial_sum_in(reg_psum_24_53), .reg_activation(reg_activation_25_53), .reg_weight(reg_weight_25_53), .reg_partial_sum(reg_psum_25_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_54( .activation_in(reg_activation_25_53), .weight_in(reg_weight_24_54), .partial_sum_in(reg_psum_24_54), .reg_activation(reg_activation_25_54), .reg_weight(reg_weight_25_54), .reg_partial_sum(reg_psum_25_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_55( .activation_in(reg_activation_25_54), .weight_in(reg_weight_24_55), .partial_sum_in(reg_psum_24_55), .reg_activation(reg_activation_25_55), .reg_weight(reg_weight_25_55), .reg_partial_sum(reg_psum_25_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_56( .activation_in(reg_activation_25_55), .weight_in(reg_weight_24_56), .partial_sum_in(reg_psum_24_56), .reg_activation(reg_activation_25_56), .reg_weight(reg_weight_25_56), .reg_partial_sum(reg_psum_25_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_57( .activation_in(reg_activation_25_56), .weight_in(reg_weight_24_57), .partial_sum_in(reg_psum_24_57), .reg_activation(reg_activation_25_57), .reg_weight(reg_weight_25_57), .reg_partial_sum(reg_psum_25_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_58( .activation_in(reg_activation_25_57), .weight_in(reg_weight_24_58), .partial_sum_in(reg_psum_24_58), .reg_activation(reg_activation_25_58), .reg_weight(reg_weight_25_58), .reg_partial_sum(reg_psum_25_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_59( .activation_in(reg_activation_25_58), .weight_in(reg_weight_24_59), .partial_sum_in(reg_psum_24_59), .reg_activation(reg_activation_25_59), .reg_weight(reg_weight_25_59), .reg_partial_sum(reg_psum_25_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_60( .activation_in(reg_activation_25_59), .weight_in(reg_weight_24_60), .partial_sum_in(reg_psum_24_60), .reg_activation(reg_activation_25_60), .reg_weight(reg_weight_25_60), .reg_partial_sum(reg_psum_25_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_61( .activation_in(reg_activation_25_60), .weight_in(reg_weight_24_61), .partial_sum_in(reg_psum_24_61), .reg_activation(reg_activation_25_61), .reg_weight(reg_weight_25_61), .reg_partial_sum(reg_psum_25_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_62( .activation_in(reg_activation_25_61), .weight_in(reg_weight_24_62), .partial_sum_in(reg_psum_24_62), .reg_activation(reg_activation_25_62), .reg_weight(reg_weight_25_62), .reg_partial_sum(reg_psum_25_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_63( .activation_in(reg_activation_25_62), .weight_in(reg_weight_24_63), .partial_sum_in(reg_psum_24_63), .reg_weight(reg_weight_25_63), .reg_partial_sum(reg_psum_25_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_0( .activation_in(in_activation_26), .weight_in(reg_weight_25_0), .partial_sum_in(reg_psum_25_0), .reg_activation(reg_activation_26_0), .reg_weight(reg_weight_26_0), .reg_partial_sum(reg_psum_26_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_1( .activation_in(reg_activation_26_0), .weight_in(reg_weight_25_1), .partial_sum_in(reg_psum_25_1), .reg_activation(reg_activation_26_1), .reg_weight(reg_weight_26_1), .reg_partial_sum(reg_psum_26_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_2( .activation_in(reg_activation_26_1), .weight_in(reg_weight_25_2), .partial_sum_in(reg_psum_25_2), .reg_activation(reg_activation_26_2), .reg_weight(reg_weight_26_2), .reg_partial_sum(reg_psum_26_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_3( .activation_in(reg_activation_26_2), .weight_in(reg_weight_25_3), .partial_sum_in(reg_psum_25_3), .reg_activation(reg_activation_26_3), .reg_weight(reg_weight_26_3), .reg_partial_sum(reg_psum_26_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_4( .activation_in(reg_activation_26_3), .weight_in(reg_weight_25_4), .partial_sum_in(reg_psum_25_4), .reg_activation(reg_activation_26_4), .reg_weight(reg_weight_26_4), .reg_partial_sum(reg_psum_26_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_5( .activation_in(reg_activation_26_4), .weight_in(reg_weight_25_5), .partial_sum_in(reg_psum_25_5), .reg_activation(reg_activation_26_5), .reg_weight(reg_weight_26_5), .reg_partial_sum(reg_psum_26_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_6( .activation_in(reg_activation_26_5), .weight_in(reg_weight_25_6), .partial_sum_in(reg_psum_25_6), .reg_activation(reg_activation_26_6), .reg_weight(reg_weight_26_6), .reg_partial_sum(reg_psum_26_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_7( .activation_in(reg_activation_26_6), .weight_in(reg_weight_25_7), .partial_sum_in(reg_psum_25_7), .reg_activation(reg_activation_26_7), .reg_weight(reg_weight_26_7), .reg_partial_sum(reg_psum_26_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_8( .activation_in(reg_activation_26_7), .weight_in(reg_weight_25_8), .partial_sum_in(reg_psum_25_8), .reg_activation(reg_activation_26_8), .reg_weight(reg_weight_26_8), .reg_partial_sum(reg_psum_26_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_9( .activation_in(reg_activation_26_8), .weight_in(reg_weight_25_9), .partial_sum_in(reg_psum_25_9), .reg_activation(reg_activation_26_9), .reg_weight(reg_weight_26_9), .reg_partial_sum(reg_psum_26_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_10( .activation_in(reg_activation_26_9), .weight_in(reg_weight_25_10), .partial_sum_in(reg_psum_25_10), .reg_activation(reg_activation_26_10), .reg_weight(reg_weight_26_10), .reg_partial_sum(reg_psum_26_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_11( .activation_in(reg_activation_26_10), .weight_in(reg_weight_25_11), .partial_sum_in(reg_psum_25_11), .reg_activation(reg_activation_26_11), .reg_weight(reg_weight_26_11), .reg_partial_sum(reg_psum_26_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_12( .activation_in(reg_activation_26_11), .weight_in(reg_weight_25_12), .partial_sum_in(reg_psum_25_12), .reg_activation(reg_activation_26_12), .reg_weight(reg_weight_26_12), .reg_partial_sum(reg_psum_26_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_13( .activation_in(reg_activation_26_12), .weight_in(reg_weight_25_13), .partial_sum_in(reg_psum_25_13), .reg_activation(reg_activation_26_13), .reg_weight(reg_weight_26_13), .reg_partial_sum(reg_psum_26_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_14( .activation_in(reg_activation_26_13), .weight_in(reg_weight_25_14), .partial_sum_in(reg_psum_25_14), .reg_activation(reg_activation_26_14), .reg_weight(reg_weight_26_14), .reg_partial_sum(reg_psum_26_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_15( .activation_in(reg_activation_26_14), .weight_in(reg_weight_25_15), .partial_sum_in(reg_psum_25_15), .reg_activation(reg_activation_26_15), .reg_weight(reg_weight_26_15), .reg_partial_sum(reg_psum_26_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_16( .activation_in(reg_activation_26_15), .weight_in(reg_weight_25_16), .partial_sum_in(reg_psum_25_16), .reg_activation(reg_activation_26_16), .reg_weight(reg_weight_26_16), .reg_partial_sum(reg_psum_26_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_17( .activation_in(reg_activation_26_16), .weight_in(reg_weight_25_17), .partial_sum_in(reg_psum_25_17), .reg_activation(reg_activation_26_17), .reg_weight(reg_weight_26_17), .reg_partial_sum(reg_psum_26_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_18( .activation_in(reg_activation_26_17), .weight_in(reg_weight_25_18), .partial_sum_in(reg_psum_25_18), .reg_activation(reg_activation_26_18), .reg_weight(reg_weight_26_18), .reg_partial_sum(reg_psum_26_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_19( .activation_in(reg_activation_26_18), .weight_in(reg_weight_25_19), .partial_sum_in(reg_psum_25_19), .reg_activation(reg_activation_26_19), .reg_weight(reg_weight_26_19), .reg_partial_sum(reg_psum_26_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_20( .activation_in(reg_activation_26_19), .weight_in(reg_weight_25_20), .partial_sum_in(reg_psum_25_20), .reg_activation(reg_activation_26_20), .reg_weight(reg_weight_26_20), .reg_partial_sum(reg_psum_26_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_21( .activation_in(reg_activation_26_20), .weight_in(reg_weight_25_21), .partial_sum_in(reg_psum_25_21), .reg_activation(reg_activation_26_21), .reg_weight(reg_weight_26_21), .reg_partial_sum(reg_psum_26_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_22( .activation_in(reg_activation_26_21), .weight_in(reg_weight_25_22), .partial_sum_in(reg_psum_25_22), .reg_activation(reg_activation_26_22), .reg_weight(reg_weight_26_22), .reg_partial_sum(reg_psum_26_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_23( .activation_in(reg_activation_26_22), .weight_in(reg_weight_25_23), .partial_sum_in(reg_psum_25_23), .reg_activation(reg_activation_26_23), .reg_weight(reg_weight_26_23), .reg_partial_sum(reg_psum_26_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_24( .activation_in(reg_activation_26_23), .weight_in(reg_weight_25_24), .partial_sum_in(reg_psum_25_24), .reg_activation(reg_activation_26_24), .reg_weight(reg_weight_26_24), .reg_partial_sum(reg_psum_26_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_25( .activation_in(reg_activation_26_24), .weight_in(reg_weight_25_25), .partial_sum_in(reg_psum_25_25), .reg_activation(reg_activation_26_25), .reg_weight(reg_weight_26_25), .reg_partial_sum(reg_psum_26_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_26( .activation_in(reg_activation_26_25), .weight_in(reg_weight_25_26), .partial_sum_in(reg_psum_25_26), .reg_activation(reg_activation_26_26), .reg_weight(reg_weight_26_26), .reg_partial_sum(reg_psum_26_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_27( .activation_in(reg_activation_26_26), .weight_in(reg_weight_25_27), .partial_sum_in(reg_psum_25_27), .reg_activation(reg_activation_26_27), .reg_weight(reg_weight_26_27), .reg_partial_sum(reg_psum_26_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_28( .activation_in(reg_activation_26_27), .weight_in(reg_weight_25_28), .partial_sum_in(reg_psum_25_28), .reg_activation(reg_activation_26_28), .reg_weight(reg_weight_26_28), .reg_partial_sum(reg_psum_26_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_29( .activation_in(reg_activation_26_28), .weight_in(reg_weight_25_29), .partial_sum_in(reg_psum_25_29), .reg_activation(reg_activation_26_29), .reg_weight(reg_weight_26_29), .reg_partial_sum(reg_psum_26_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_30( .activation_in(reg_activation_26_29), .weight_in(reg_weight_25_30), .partial_sum_in(reg_psum_25_30), .reg_activation(reg_activation_26_30), .reg_weight(reg_weight_26_30), .reg_partial_sum(reg_psum_26_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_31( .activation_in(reg_activation_26_30), .weight_in(reg_weight_25_31), .partial_sum_in(reg_psum_25_31), .reg_activation(reg_activation_26_31), .reg_weight(reg_weight_26_31), .reg_partial_sum(reg_psum_26_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_32( .activation_in(reg_activation_26_31), .weight_in(reg_weight_25_32), .partial_sum_in(reg_psum_25_32), .reg_activation(reg_activation_26_32), .reg_weight(reg_weight_26_32), .reg_partial_sum(reg_psum_26_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_33( .activation_in(reg_activation_26_32), .weight_in(reg_weight_25_33), .partial_sum_in(reg_psum_25_33), .reg_activation(reg_activation_26_33), .reg_weight(reg_weight_26_33), .reg_partial_sum(reg_psum_26_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_34( .activation_in(reg_activation_26_33), .weight_in(reg_weight_25_34), .partial_sum_in(reg_psum_25_34), .reg_activation(reg_activation_26_34), .reg_weight(reg_weight_26_34), .reg_partial_sum(reg_psum_26_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_35( .activation_in(reg_activation_26_34), .weight_in(reg_weight_25_35), .partial_sum_in(reg_psum_25_35), .reg_activation(reg_activation_26_35), .reg_weight(reg_weight_26_35), .reg_partial_sum(reg_psum_26_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_36( .activation_in(reg_activation_26_35), .weight_in(reg_weight_25_36), .partial_sum_in(reg_psum_25_36), .reg_activation(reg_activation_26_36), .reg_weight(reg_weight_26_36), .reg_partial_sum(reg_psum_26_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_37( .activation_in(reg_activation_26_36), .weight_in(reg_weight_25_37), .partial_sum_in(reg_psum_25_37), .reg_activation(reg_activation_26_37), .reg_weight(reg_weight_26_37), .reg_partial_sum(reg_psum_26_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_38( .activation_in(reg_activation_26_37), .weight_in(reg_weight_25_38), .partial_sum_in(reg_psum_25_38), .reg_activation(reg_activation_26_38), .reg_weight(reg_weight_26_38), .reg_partial_sum(reg_psum_26_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_39( .activation_in(reg_activation_26_38), .weight_in(reg_weight_25_39), .partial_sum_in(reg_psum_25_39), .reg_activation(reg_activation_26_39), .reg_weight(reg_weight_26_39), .reg_partial_sum(reg_psum_26_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_40( .activation_in(reg_activation_26_39), .weight_in(reg_weight_25_40), .partial_sum_in(reg_psum_25_40), .reg_activation(reg_activation_26_40), .reg_weight(reg_weight_26_40), .reg_partial_sum(reg_psum_26_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_41( .activation_in(reg_activation_26_40), .weight_in(reg_weight_25_41), .partial_sum_in(reg_psum_25_41), .reg_activation(reg_activation_26_41), .reg_weight(reg_weight_26_41), .reg_partial_sum(reg_psum_26_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_42( .activation_in(reg_activation_26_41), .weight_in(reg_weight_25_42), .partial_sum_in(reg_psum_25_42), .reg_activation(reg_activation_26_42), .reg_weight(reg_weight_26_42), .reg_partial_sum(reg_psum_26_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_43( .activation_in(reg_activation_26_42), .weight_in(reg_weight_25_43), .partial_sum_in(reg_psum_25_43), .reg_activation(reg_activation_26_43), .reg_weight(reg_weight_26_43), .reg_partial_sum(reg_psum_26_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_44( .activation_in(reg_activation_26_43), .weight_in(reg_weight_25_44), .partial_sum_in(reg_psum_25_44), .reg_activation(reg_activation_26_44), .reg_weight(reg_weight_26_44), .reg_partial_sum(reg_psum_26_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_45( .activation_in(reg_activation_26_44), .weight_in(reg_weight_25_45), .partial_sum_in(reg_psum_25_45), .reg_activation(reg_activation_26_45), .reg_weight(reg_weight_26_45), .reg_partial_sum(reg_psum_26_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_46( .activation_in(reg_activation_26_45), .weight_in(reg_weight_25_46), .partial_sum_in(reg_psum_25_46), .reg_activation(reg_activation_26_46), .reg_weight(reg_weight_26_46), .reg_partial_sum(reg_psum_26_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_47( .activation_in(reg_activation_26_46), .weight_in(reg_weight_25_47), .partial_sum_in(reg_psum_25_47), .reg_activation(reg_activation_26_47), .reg_weight(reg_weight_26_47), .reg_partial_sum(reg_psum_26_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_48( .activation_in(reg_activation_26_47), .weight_in(reg_weight_25_48), .partial_sum_in(reg_psum_25_48), .reg_activation(reg_activation_26_48), .reg_weight(reg_weight_26_48), .reg_partial_sum(reg_psum_26_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_49( .activation_in(reg_activation_26_48), .weight_in(reg_weight_25_49), .partial_sum_in(reg_psum_25_49), .reg_activation(reg_activation_26_49), .reg_weight(reg_weight_26_49), .reg_partial_sum(reg_psum_26_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_50( .activation_in(reg_activation_26_49), .weight_in(reg_weight_25_50), .partial_sum_in(reg_psum_25_50), .reg_activation(reg_activation_26_50), .reg_weight(reg_weight_26_50), .reg_partial_sum(reg_psum_26_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_51( .activation_in(reg_activation_26_50), .weight_in(reg_weight_25_51), .partial_sum_in(reg_psum_25_51), .reg_activation(reg_activation_26_51), .reg_weight(reg_weight_26_51), .reg_partial_sum(reg_psum_26_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_52( .activation_in(reg_activation_26_51), .weight_in(reg_weight_25_52), .partial_sum_in(reg_psum_25_52), .reg_activation(reg_activation_26_52), .reg_weight(reg_weight_26_52), .reg_partial_sum(reg_psum_26_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_53( .activation_in(reg_activation_26_52), .weight_in(reg_weight_25_53), .partial_sum_in(reg_psum_25_53), .reg_activation(reg_activation_26_53), .reg_weight(reg_weight_26_53), .reg_partial_sum(reg_psum_26_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_54( .activation_in(reg_activation_26_53), .weight_in(reg_weight_25_54), .partial_sum_in(reg_psum_25_54), .reg_activation(reg_activation_26_54), .reg_weight(reg_weight_26_54), .reg_partial_sum(reg_psum_26_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_55( .activation_in(reg_activation_26_54), .weight_in(reg_weight_25_55), .partial_sum_in(reg_psum_25_55), .reg_activation(reg_activation_26_55), .reg_weight(reg_weight_26_55), .reg_partial_sum(reg_psum_26_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_56( .activation_in(reg_activation_26_55), .weight_in(reg_weight_25_56), .partial_sum_in(reg_psum_25_56), .reg_activation(reg_activation_26_56), .reg_weight(reg_weight_26_56), .reg_partial_sum(reg_psum_26_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_57( .activation_in(reg_activation_26_56), .weight_in(reg_weight_25_57), .partial_sum_in(reg_psum_25_57), .reg_activation(reg_activation_26_57), .reg_weight(reg_weight_26_57), .reg_partial_sum(reg_psum_26_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_58( .activation_in(reg_activation_26_57), .weight_in(reg_weight_25_58), .partial_sum_in(reg_psum_25_58), .reg_activation(reg_activation_26_58), .reg_weight(reg_weight_26_58), .reg_partial_sum(reg_psum_26_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_59( .activation_in(reg_activation_26_58), .weight_in(reg_weight_25_59), .partial_sum_in(reg_psum_25_59), .reg_activation(reg_activation_26_59), .reg_weight(reg_weight_26_59), .reg_partial_sum(reg_psum_26_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_60( .activation_in(reg_activation_26_59), .weight_in(reg_weight_25_60), .partial_sum_in(reg_psum_25_60), .reg_activation(reg_activation_26_60), .reg_weight(reg_weight_26_60), .reg_partial_sum(reg_psum_26_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_61( .activation_in(reg_activation_26_60), .weight_in(reg_weight_25_61), .partial_sum_in(reg_psum_25_61), .reg_activation(reg_activation_26_61), .reg_weight(reg_weight_26_61), .reg_partial_sum(reg_psum_26_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_62( .activation_in(reg_activation_26_61), .weight_in(reg_weight_25_62), .partial_sum_in(reg_psum_25_62), .reg_activation(reg_activation_26_62), .reg_weight(reg_weight_26_62), .reg_partial_sum(reg_psum_26_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_63( .activation_in(reg_activation_26_62), .weight_in(reg_weight_25_63), .partial_sum_in(reg_psum_25_63), .reg_weight(reg_weight_26_63), .reg_partial_sum(reg_psum_26_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_0( .activation_in(in_activation_27), .weight_in(reg_weight_26_0), .partial_sum_in(reg_psum_26_0), .reg_activation(reg_activation_27_0), .reg_weight(reg_weight_27_0), .reg_partial_sum(reg_psum_27_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_1( .activation_in(reg_activation_27_0), .weight_in(reg_weight_26_1), .partial_sum_in(reg_psum_26_1), .reg_activation(reg_activation_27_1), .reg_weight(reg_weight_27_1), .reg_partial_sum(reg_psum_27_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_2( .activation_in(reg_activation_27_1), .weight_in(reg_weight_26_2), .partial_sum_in(reg_psum_26_2), .reg_activation(reg_activation_27_2), .reg_weight(reg_weight_27_2), .reg_partial_sum(reg_psum_27_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_3( .activation_in(reg_activation_27_2), .weight_in(reg_weight_26_3), .partial_sum_in(reg_psum_26_3), .reg_activation(reg_activation_27_3), .reg_weight(reg_weight_27_3), .reg_partial_sum(reg_psum_27_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_4( .activation_in(reg_activation_27_3), .weight_in(reg_weight_26_4), .partial_sum_in(reg_psum_26_4), .reg_activation(reg_activation_27_4), .reg_weight(reg_weight_27_4), .reg_partial_sum(reg_psum_27_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_5( .activation_in(reg_activation_27_4), .weight_in(reg_weight_26_5), .partial_sum_in(reg_psum_26_5), .reg_activation(reg_activation_27_5), .reg_weight(reg_weight_27_5), .reg_partial_sum(reg_psum_27_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_6( .activation_in(reg_activation_27_5), .weight_in(reg_weight_26_6), .partial_sum_in(reg_psum_26_6), .reg_activation(reg_activation_27_6), .reg_weight(reg_weight_27_6), .reg_partial_sum(reg_psum_27_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_7( .activation_in(reg_activation_27_6), .weight_in(reg_weight_26_7), .partial_sum_in(reg_psum_26_7), .reg_activation(reg_activation_27_7), .reg_weight(reg_weight_27_7), .reg_partial_sum(reg_psum_27_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_8( .activation_in(reg_activation_27_7), .weight_in(reg_weight_26_8), .partial_sum_in(reg_psum_26_8), .reg_activation(reg_activation_27_8), .reg_weight(reg_weight_27_8), .reg_partial_sum(reg_psum_27_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_9( .activation_in(reg_activation_27_8), .weight_in(reg_weight_26_9), .partial_sum_in(reg_psum_26_9), .reg_activation(reg_activation_27_9), .reg_weight(reg_weight_27_9), .reg_partial_sum(reg_psum_27_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_10( .activation_in(reg_activation_27_9), .weight_in(reg_weight_26_10), .partial_sum_in(reg_psum_26_10), .reg_activation(reg_activation_27_10), .reg_weight(reg_weight_27_10), .reg_partial_sum(reg_psum_27_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_11( .activation_in(reg_activation_27_10), .weight_in(reg_weight_26_11), .partial_sum_in(reg_psum_26_11), .reg_activation(reg_activation_27_11), .reg_weight(reg_weight_27_11), .reg_partial_sum(reg_psum_27_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_12( .activation_in(reg_activation_27_11), .weight_in(reg_weight_26_12), .partial_sum_in(reg_psum_26_12), .reg_activation(reg_activation_27_12), .reg_weight(reg_weight_27_12), .reg_partial_sum(reg_psum_27_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_13( .activation_in(reg_activation_27_12), .weight_in(reg_weight_26_13), .partial_sum_in(reg_psum_26_13), .reg_activation(reg_activation_27_13), .reg_weight(reg_weight_27_13), .reg_partial_sum(reg_psum_27_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_14( .activation_in(reg_activation_27_13), .weight_in(reg_weight_26_14), .partial_sum_in(reg_psum_26_14), .reg_activation(reg_activation_27_14), .reg_weight(reg_weight_27_14), .reg_partial_sum(reg_psum_27_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_15( .activation_in(reg_activation_27_14), .weight_in(reg_weight_26_15), .partial_sum_in(reg_psum_26_15), .reg_activation(reg_activation_27_15), .reg_weight(reg_weight_27_15), .reg_partial_sum(reg_psum_27_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_16( .activation_in(reg_activation_27_15), .weight_in(reg_weight_26_16), .partial_sum_in(reg_psum_26_16), .reg_activation(reg_activation_27_16), .reg_weight(reg_weight_27_16), .reg_partial_sum(reg_psum_27_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_17( .activation_in(reg_activation_27_16), .weight_in(reg_weight_26_17), .partial_sum_in(reg_psum_26_17), .reg_activation(reg_activation_27_17), .reg_weight(reg_weight_27_17), .reg_partial_sum(reg_psum_27_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_18( .activation_in(reg_activation_27_17), .weight_in(reg_weight_26_18), .partial_sum_in(reg_psum_26_18), .reg_activation(reg_activation_27_18), .reg_weight(reg_weight_27_18), .reg_partial_sum(reg_psum_27_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_19( .activation_in(reg_activation_27_18), .weight_in(reg_weight_26_19), .partial_sum_in(reg_psum_26_19), .reg_activation(reg_activation_27_19), .reg_weight(reg_weight_27_19), .reg_partial_sum(reg_psum_27_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_20( .activation_in(reg_activation_27_19), .weight_in(reg_weight_26_20), .partial_sum_in(reg_psum_26_20), .reg_activation(reg_activation_27_20), .reg_weight(reg_weight_27_20), .reg_partial_sum(reg_psum_27_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_21( .activation_in(reg_activation_27_20), .weight_in(reg_weight_26_21), .partial_sum_in(reg_psum_26_21), .reg_activation(reg_activation_27_21), .reg_weight(reg_weight_27_21), .reg_partial_sum(reg_psum_27_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_22( .activation_in(reg_activation_27_21), .weight_in(reg_weight_26_22), .partial_sum_in(reg_psum_26_22), .reg_activation(reg_activation_27_22), .reg_weight(reg_weight_27_22), .reg_partial_sum(reg_psum_27_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_23( .activation_in(reg_activation_27_22), .weight_in(reg_weight_26_23), .partial_sum_in(reg_psum_26_23), .reg_activation(reg_activation_27_23), .reg_weight(reg_weight_27_23), .reg_partial_sum(reg_psum_27_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_24( .activation_in(reg_activation_27_23), .weight_in(reg_weight_26_24), .partial_sum_in(reg_psum_26_24), .reg_activation(reg_activation_27_24), .reg_weight(reg_weight_27_24), .reg_partial_sum(reg_psum_27_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_25( .activation_in(reg_activation_27_24), .weight_in(reg_weight_26_25), .partial_sum_in(reg_psum_26_25), .reg_activation(reg_activation_27_25), .reg_weight(reg_weight_27_25), .reg_partial_sum(reg_psum_27_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_26( .activation_in(reg_activation_27_25), .weight_in(reg_weight_26_26), .partial_sum_in(reg_psum_26_26), .reg_activation(reg_activation_27_26), .reg_weight(reg_weight_27_26), .reg_partial_sum(reg_psum_27_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_27( .activation_in(reg_activation_27_26), .weight_in(reg_weight_26_27), .partial_sum_in(reg_psum_26_27), .reg_activation(reg_activation_27_27), .reg_weight(reg_weight_27_27), .reg_partial_sum(reg_psum_27_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_28( .activation_in(reg_activation_27_27), .weight_in(reg_weight_26_28), .partial_sum_in(reg_psum_26_28), .reg_activation(reg_activation_27_28), .reg_weight(reg_weight_27_28), .reg_partial_sum(reg_psum_27_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_29( .activation_in(reg_activation_27_28), .weight_in(reg_weight_26_29), .partial_sum_in(reg_psum_26_29), .reg_activation(reg_activation_27_29), .reg_weight(reg_weight_27_29), .reg_partial_sum(reg_psum_27_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_30( .activation_in(reg_activation_27_29), .weight_in(reg_weight_26_30), .partial_sum_in(reg_psum_26_30), .reg_activation(reg_activation_27_30), .reg_weight(reg_weight_27_30), .reg_partial_sum(reg_psum_27_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_31( .activation_in(reg_activation_27_30), .weight_in(reg_weight_26_31), .partial_sum_in(reg_psum_26_31), .reg_activation(reg_activation_27_31), .reg_weight(reg_weight_27_31), .reg_partial_sum(reg_psum_27_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_32( .activation_in(reg_activation_27_31), .weight_in(reg_weight_26_32), .partial_sum_in(reg_psum_26_32), .reg_activation(reg_activation_27_32), .reg_weight(reg_weight_27_32), .reg_partial_sum(reg_psum_27_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_33( .activation_in(reg_activation_27_32), .weight_in(reg_weight_26_33), .partial_sum_in(reg_psum_26_33), .reg_activation(reg_activation_27_33), .reg_weight(reg_weight_27_33), .reg_partial_sum(reg_psum_27_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_34( .activation_in(reg_activation_27_33), .weight_in(reg_weight_26_34), .partial_sum_in(reg_psum_26_34), .reg_activation(reg_activation_27_34), .reg_weight(reg_weight_27_34), .reg_partial_sum(reg_psum_27_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_35( .activation_in(reg_activation_27_34), .weight_in(reg_weight_26_35), .partial_sum_in(reg_psum_26_35), .reg_activation(reg_activation_27_35), .reg_weight(reg_weight_27_35), .reg_partial_sum(reg_psum_27_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_36( .activation_in(reg_activation_27_35), .weight_in(reg_weight_26_36), .partial_sum_in(reg_psum_26_36), .reg_activation(reg_activation_27_36), .reg_weight(reg_weight_27_36), .reg_partial_sum(reg_psum_27_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_37( .activation_in(reg_activation_27_36), .weight_in(reg_weight_26_37), .partial_sum_in(reg_psum_26_37), .reg_activation(reg_activation_27_37), .reg_weight(reg_weight_27_37), .reg_partial_sum(reg_psum_27_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_38( .activation_in(reg_activation_27_37), .weight_in(reg_weight_26_38), .partial_sum_in(reg_psum_26_38), .reg_activation(reg_activation_27_38), .reg_weight(reg_weight_27_38), .reg_partial_sum(reg_psum_27_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_39( .activation_in(reg_activation_27_38), .weight_in(reg_weight_26_39), .partial_sum_in(reg_psum_26_39), .reg_activation(reg_activation_27_39), .reg_weight(reg_weight_27_39), .reg_partial_sum(reg_psum_27_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_40( .activation_in(reg_activation_27_39), .weight_in(reg_weight_26_40), .partial_sum_in(reg_psum_26_40), .reg_activation(reg_activation_27_40), .reg_weight(reg_weight_27_40), .reg_partial_sum(reg_psum_27_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_41( .activation_in(reg_activation_27_40), .weight_in(reg_weight_26_41), .partial_sum_in(reg_psum_26_41), .reg_activation(reg_activation_27_41), .reg_weight(reg_weight_27_41), .reg_partial_sum(reg_psum_27_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_42( .activation_in(reg_activation_27_41), .weight_in(reg_weight_26_42), .partial_sum_in(reg_psum_26_42), .reg_activation(reg_activation_27_42), .reg_weight(reg_weight_27_42), .reg_partial_sum(reg_psum_27_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_43( .activation_in(reg_activation_27_42), .weight_in(reg_weight_26_43), .partial_sum_in(reg_psum_26_43), .reg_activation(reg_activation_27_43), .reg_weight(reg_weight_27_43), .reg_partial_sum(reg_psum_27_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_44( .activation_in(reg_activation_27_43), .weight_in(reg_weight_26_44), .partial_sum_in(reg_psum_26_44), .reg_activation(reg_activation_27_44), .reg_weight(reg_weight_27_44), .reg_partial_sum(reg_psum_27_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_45( .activation_in(reg_activation_27_44), .weight_in(reg_weight_26_45), .partial_sum_in(reg_psum_26_45), .reg_activation(reg_activation_27_45), .reg_weight(reg_weight_27_45), .reg_partial_sum(reg_psum_27_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_46( .activation_in(reg_activation_27_45), .weight_in(reg_weight_26_46), .partial_sum_in(reg_psum_26_46), .reg_activation(reg_activation_27_46), .reg_weight(reg_weight_27_46), .reg_partial_sum(reg_psum_27_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_47( .activation_in(reg_activation_27_46), .weight_in(reg_weight_26_47), .partial_sum_in(reg_psum_26_47), .reg_activation(reg_activation_27_47), .reg_weight(reg_weight_27_47), .reg_partial_sum(reg_psum_27_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_48( .activation_in(reg_activation_27_47), .weight_in(reg_weight_26_48), .partial_sum_in(reg_psum_26_48), .reg_activation(reg_activation_27_48), .reg_weight(reg_weight_27_48), .reg_partial_sum(reg_psum_27_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_49( .activation_in(reg_activation_27_48), .weight_in(reg_weight_26_49), .partial_sum_in(reg_psum_26_49), .reg_activation(reg_activation_27_49), .reg_weight(reg_weight_27_49), .reg_partial_sum(reg_psum_27_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_50( .activation_in(reg_activation_27_49), .weight_in(reg_weight_26_50), .partial_sum_in(reg_psum_26_50), .reg_activation(reg_activation_27_50), .reg_weight(reg_weight_27_50), .reg_partial_sum(reg_psum_27_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_51( .activation_in(reg_activation_27_50), .weight_in(reg_weight_26_51), .partial_sum_in(reg_psum_26_51), .reg_activation(reg_activation_27_51), .reg_weight(reg_weight_27_51), .reg_partial_sum(reg_psum_27_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_52( .activation_in(reg_activation_27_51), .weight_in(reg_weight_26_52), .partial_sum_in(reg_psum_26_52), .reg_activation(reg_activation_27_52), .reg_weight(reg_weight_27_52), .reg_partial_sum(reg_psum_27_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_53( .activation_in(reg_activation_27_52), .weight_in(reg_weight_26_53), .partial_sum_in(reg_psum_26_53), .reg_activation(reg_activation_27_53), .reg_weight(reg_weight_27_53), .reg_partial_sum(reg_psum_27_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_54( .activation_in(reg_activation_27_53), .weight_in(reg_weight_26_54), .partial_sum_in(reg_psum_26_54), .reg_activation(reg_activation_27_54), .reg_weight(reg_weight_27_54), .reg_partial_sum(reg_psum_27_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_55( .activation_in(reg_activation_27_54), .weight_in(reg_weight_26_55), .partial_sum_in(reg_psum_26_55), .reg_activation(reg_activation_27_55), .reg_weight(reg_weight_27_55), .reg_partial_sum(reg_psum_27_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_56( .activation_in(reg_activation_27_55), .weight_in(reg_weight_26_56), .partial_sum_in(reg_psum_26_56), .reg_activation(reg_activation_27_56), .reg_weight(reg_weight_27_56), .reg_partial_sum(reg_psum_27_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_57( .activation_in(reg_activation_27_56), .weight_in(reg_weight_26_57), .partial_sum_in(reg_psum_26_57), .reg_activation(reg_activation_27_57), .reg_weight(reg_weight_27_57), .reg_partial_sum(reg_psum_27_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_58( .activation_in(reg_activation_27_57), .weight_in(reg_weight_26_58), .partial_sum_in(reg_psum_26_58), .reg_activation(reg_activation_27_58), .reg_weight(reg_weight_27_58), .reg_partial_sum(reg_psum_27_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_59( .activation_in(reg_activation_27_58), .weight_in(reg_weight_26_59), .partial_sum_in(reg_psum_26_59), .reg_activation(reg_activation_27_59), .reg_weight(reg_weight_27_59), .reg_partial_sum(reg_psum_27_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_60( .activation_in(reg_activation_27_59), .weight_in(reg_weight_26_60), .partial_sum_in(reg_psum_26_60), .reg_activation(reg_activation_27_60), .reg_weight(reg_weight_27_60), .reg_partial_sum(reg_psum_27_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_61( .activation_in(reg_activation_27_60), .weight_in(reg_weight_26_61), .partial_sum_in(reg_psum_26_61), .reg_activation(reg_activation_27_61), .reg_weight(reg_weight_27_61), .reg_partial_sum(reg_psum_27_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_62( .activation_in(reg_activation_27_61), .weight_in(reg_weight_26_62), .partial_sum_in(reg_psum_26_62), .reg_activation(reg_activation_27_62), .reg_weight(reg_weight_27_62), .reg_partial_sum(reg_psum_27_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_63( .activation_in(reg_activation_27_62), .weight_in(reg_weight_26_63), .partial_sum_in(reg_psum_26_63), .reg_weight(reg_weight_27_63), .reg_partial_sum(reg_psum_27_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_0( .activation_in(in_activation_28), .weight_in(reg_weight_27_0), .partial_sum_in(reg_psum_27_0), .reg_activation(reg_activation_28_0), .reg_weight(reg_weight_28_0), .reg_partial_sum(reg_psum_28_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_1( .activation_in(reg_activation_28_0), .weight_in(reg_weight_27_1), .partial_sum_in(reg_psum_27_1), .reg_activation(reg_activation_28_1), .reg_weight(reg_weight_28_1), .reg_partial_sum(reg_psum_28_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_2( .activation_in(reg_activation_28_1), .weight_in(reg_weight_27_2), .partial_sum_in(reg_psum_27_2), .reg_activation(reg_activation_28_2), .reg_weight(reg_weight_28_2), .reg_partial_sum(reg_psum_28_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_3( .activation_in(reg_activation_28_2), .weight_in(reg_weight_27_3), .partial_sum_in(reg_psum_27_3), .reg_activation(reg_activation_28_3), .reg_weight(reg_weight_28_3), .reg_partial_sum(reg_psum_28_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_4( .activation_in(reg_activation_28_3), .weight_in(reg_weight_27_4), .partial_sum_in(reg_psum_27_4), .reg_activation(reg_activation_28_4), .reg_weight(reg_weight_28_4), .reg_partial_sum(reg_psum_28_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_5( .activation_in(reg_activation_28_4), .weight_in(reg_weight_27_5), .partial_sum_in(reg_psum_27_5), .reg_activation(reg_activation_28_5), .reg_weight(reg_weight_28_5), .reg_partial_sum(reg_psum_28_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_6( .activation_in(reg_activation_28_5), .weight_in(reg_weight_27_6), .partial_sum_in(reg_psum_27_6), .reg_activation(reg_activation_28_6), .reg_weight(reg_weight_28_6), .reg_partial_sum(reg_psum_28_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_7( .activation_in(reg_activation_28_6), .weight_in(reg_weight_27_7), .partial_sum_in(reg_psum_27_7), .reg_activation(reg_activation_28_7), .reg_weight(reg_weight_28_7), .reg_partial_sum(reg_psum_28_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_8( .activation_in(reg_activation_28_7), .weight_in(reg_weight_27_8), .partial_sum_in(reg_psum_27_8), .reg_activation(reg_activation_28_8), .reg_weight(reg_weight_28_8), .reg_partial_sum(reg_psum_28_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_9( .activation_in(reg_activation_28_8), .weight_in(reg_weight_27_9), .partial_sum_in(reg_psum_27_9), .reg_activation(reg_activation_28_9), .reg_weight(reg_weight_28_9), .reg_partial_sum(reg_psum_28_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_10( .activation_in(reg_activation_28_9), .weight_in(reg_weight_27_10), .partial_sum_in(reg_psum_27_10), .reg_activation(reg_activation_28_10), .reg_weight(reg_weight_28_10), .reg_partial_sum(reg_psum_28_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_11( .activation_in(reg_activation_28_10), .weight_in(reg_weight_27_11), .partial_sum_in(reg_psum_27_11), .reg_activation(reg_activation_28_11), .reg_weight(reg_weight_28_11), .reg_partial_sum(reg_psum_28_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_12( .activation_in(reg_activation_28_11), .weight_in(reg_weight_27_12), .partial_sum_in(reg_psum_27_12), .reg_activation(reg_activation_28_12), .reg_weight(reg_weight_28_12), .reg_partial_sum(reg_psum_28_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_13( .activation_in(reg_activation_28_12), .weight_in(reg_weight_27_13), .partial_sum_in(reg_psum_27_13), .reg_activation(reg_activation_28_13), .reg_weight(reg_weight_28_13), .reg_partial_sum(reg_psum_28_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_14( .activation_in(reg_activation_28_13), .weight_in(reg_weight_27_14), .partial_sum_in(reg_psum_27_14), .reg_activation(reg_activation_28_14), .reg_weight(reg_weight_28_14), .reg_partial_sum(reg_psum_28_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_15( .activation_in(reg_activation_28_14), .weight_in(reg_weight_27_15), .partial_sum_in(reg_psum_27_15), .reg_activation(reg_activation_28_15), .reg_weight(reg_weight_28_15), .reg_partial_sum(reg_psum_28_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_16( .activation_in(reg_activation_28_15), .weight_in(reg_weight_27_16), .partial_sum_in(reg_psum_27_16), .reg_activation(reg_activation_28_16), .reg_weight(reg_weight_28_16), .reg_partial_sum(reg_psum_28_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_17( .activation_in(reg_activation_28_16), .weight_in(reg_weight_27_17), .partial_sum_in(reg_psum_27_17), .reg_activation(reg_activation_28_17), .reg_weight(reg_weight_28_17), .reg_partial_sum(reg_psum_28_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_18( .activation_in(reg_activation_28_17), .weight_in(reg_weight_27_18), .partial_sum_in(reg_psum_27_18), .reg_activation(reg_activation_28_18), .reg_weight(reg_weight_28_18), .reg_partial_sum(reg_psum_28_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_19( .activation_in(reg_activation_28_18), .weight_in(reg_weight_27_19), .partial_sum_in(reg_psum_27_19), .reg_activation(reg_activation_28_19), .reg_weight(reg_weight_28_19), .reg_partial_sum(reg_psum_28_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_20( .activation_in(reg_activation_28_19), .weight_in(reg_weight_27_20), .partial_sum_in(reg_psum_27_20), .reg_activation(reg_activation_28_20), .reg_weight(reg_weight_28_20), .reg_partial_sum(reg_psum_28_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_21( .activation_in(reg_activation_28_20), .weight_in(reg_weight_27_21), .partial_sum_in(reg_psum_27_21), .reg_activation(reg_activation_28_21), .reg_weight(reg_weight_28_21), .reg_partial_sum(reg_psum_28_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_22( .activation_in(reg_activation_28_21), .weight_in(reg_weight_27_22), .partial_sum_in(reg_psum_27_22), .reg_activation(reg_activation_28_22), .reg_weight(reg_weight_28_22), .reg_partial_sum(reg_psum_28_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_23( .activation_in(reg_activation_28_22), .weight_in(reg_weight_27_23), .partial_sum_in(reg_psum_27_23), .reg_activation(reg_activation_28_23), .reg_weight(reg_weight_28_23), .reg_partial_sum(reg_psum_28_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_24( .activation_in(reg_activation_28_23), .weight_in(reg_weight_27_24), .partial_sum_in(reg_psum_27_24), .reg_activation(reg_activation_28_24), .reg_weight(reg_weight_28_24), .reg_partial_sum(reg_psum_28_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_25( .activation_in(reg_activation_28_24), .weight_in(reg_weight_27_25), .partial_sum_in(reg_psum_27_25), .reg_activation(reg_activation_28_25), .reg_weight(reg_weight_28_25), .reg_partial_sum(reg_psum_28_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_26( .activation_in(reg_activation_28_25), .weight_in(reg_weight_27_26), .partial_sum_in(reg_psum_27_26), .reg_activation(reg_activation_28_26), .reg_weight(reg_weight_28_26), .reg_partial_sum(reg_psum_28_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_27( .activation_in(reg_activation_28_26), .weight_in(reg_weight_27_27), .partial_sum_in(reg_psum_27_27), .reg_activation(reg_activation_28_27), .reg_weight(reg_weight_28_27), .reg_partial_sum(reg_psum_28_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_28( .activation_in(reg_activation_28_27), .weight_in(reg_weight_27_28), .partial_sum_in(reg_psum_27_28), .reg_activation(reg_activation_28_28), .reg_weight(reg_weight_28_28), .reg_partial_sum(reg_psum_28_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_29( .activation_in(reg_activation_28_28), .weight_in(reg_weight_27_29), .partial_sum_in(reg_psum_27_29), .reg_activation(reg_activation_28_29), .reg_weight(reg_weight_28_29), .reg_partial_sum(reg_psum_28_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_30( .activation_in(reg_activation_28_29), .weight_in(reg_weight_27_30), .partial_sum_in(reg_psum_27_30), .reg_activation(reg_activation_28_30), .reg_weight(reg_weight_28_30), .reg_partial_sum(reg_psum_28_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_31( .activation_in(reg_activation_28_30), .weight_in(reg_weight_27_31), .partial_sum_in(reg_psum_27_31), .reg_activation(reg_activation_28_31), .reg_weight(reg_weight_28_31), .reg_partial_sum(reg_psum_28_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_32( .activation_in(reg_activation_28_31), .weight_in(reg_weight_27_32), .partial_sum_in(reg_psum_27_32), .reg_activation(reg_activation_28_32), .reg_weight(reg_weight_28_32), .reg_partial_sum(reg_psum_28_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_33( .activation_in(reg_activation_28_32), .weight_in(reg_weight_27_33), .partial_sum_in(reg_psum_27_33), .reg_activation(reg_activation_28_33), .reg_weight(reg_weight_28_33), .reg_partial_sum(reg_psum_28_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_34( .activation_in(reg_activation_28_33), .weight_in(reg_weight_27_34), .partial_sum_in(reg_psum_27_34), .reg_activation(reg_activation_28_34), .reg_weight(reg_weight_28_34), .reg_partial_sum(reg_psum_28_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_35( .activation_in(reg_activation_28_34), .weight_in(reg_weight_27_35), .partial_sum_in(reg_psum_27_35), .reg_activation(reg_activation_28_35), .reg_weight(reg_weight_28_35), .reg_partial_sum(reg_psum_28_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_36( .activation_in(reg_activation_28_35), .weight_in(reg_weight_27_36), .partial_sum_in(reg_psum_27_36), .reg_activation(reg_activation_28_36), .reg_weight(reg_weight_28_36), .reg_partial_sum(reg_psum_28_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_37( .activation_in(reg_activation_28_36), .weight_in(reg_weight_27_37), .partial_sum_in(reg_psum_27_37), .reg_activation(reg_activation_28_37), .reg_weight(reg_weight_28_37), .reg_partial_sum(reg_psum_28_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_38( .activation_in(reg_activation_28_37), .weight_in(reg_weight_27_38), .partial_sum_in(reg_psum_27_38), .reg_activation(reg_activation_28_38), .reg_weight(reg_weight_28_38), .reg_partial_sum(reg_psum_28_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_39( .activation_in(reg_activation_28_38), .weight_in(reg_weight_27_39), .partial_sum_in(reg_psum_27_39), .reg_activation(reg_activation_28_39), .reg_weight(reg_weight_28_39), .reg_partial_sum(reg_psum_28_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_40( .activation_in(reg_activation_28_39), .weight_in(reg_weight_27_40), .partial_sum_in(reg_psum_27_40), .reg_activation(reg_activation_28_40), .reg_weight(reg_weight_28_40), .reg_partial_sum(reg_psum_28_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_41( .activation_in(reg_activation_28_40), .weight_in(reg_weight_27_41), .partial_sum_in(reg_psum_27_41), .reg_activation(reg_activation_28_41), .reg_weight(reg_weight_28_41), .reg_partial_sum(reg_psum_28_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_42( .activation_in(reg_activation_28_41), .weight_in(reg_weight_27_42), .partial_sum_in(reg_psum_27_42), .reg_activation(reg_activation_28_42), .reg_weight(reg_weight_28_42), .reg_partial_sum(reg_psum_28_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_43( .activation_in(reg_activation_28_42), .weight_in(reg_weight_27_43), .partial_sum_in(reg_psum_27_43), .reg_activation(reg_activation_28_43), .reg_weight(reg_weight_28_43), .reg_partial_sum(reg_psum_28_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_44( .activation_in(reg_activation_28_43), .weight_in(reg_weight_27_44), .partial_sum_in(reg_psum_27_44), .reg_activation(reg_activation_28_44), .reg_weight(reg_weight_28_44), .reg_partial_sum(reg_psum_28_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_45( .activation_in(reg_activation_28_44), .weight_in(reg_weight_27_45), .partial_sum_in(reg_psum_27_45), .reg_activation(reg_activation_28_45), .reg_weight(reg_weight_28_45), .reg_partial_sum(reg_psum_28_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_46( .activation_in(reg_activation_28_45), .weight_in(reg_weight_27_46), .partial_sum_in(reg_psum_27_46), .reg_activation(reg_activation_28_46), .reg_weight(reg_weight_28_46), .reg_partial_sum(reg_psum_28_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_47( .activation_in(reg_activation_28_46), .weight_in(reg_weight_27_47), .partial_sum_in(reg_psum_27_47), .reg_activation(reg_activation_28_47), .reg_weight(reg_weight_28_47), .reg_partial_sum(reg_psum_28_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_48( .activation_in(reg_activation_28_47), .weight_in(reg_weight_27_48), .partial_sum_in(reg_psum_27_48), .reg_activation(reg_activation_28_48), .reg_weight(reg_weight_28_48), .reg_partial_sum(reg_psum_28_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_49( .activation_in(reg_activation_28_48), .weight_in(reg_weight_27_49), .partial_sum_in(reg_psum_27_49), .reg_activation(reg_activation_28_49), .reg_weight(reg_weight_28_49), .reg_partial_sum(reg_psum_28_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_50( .activation_in(reg_activation_28_49), .weight_in(reg_weight_27_50), .partial_sum_in(reg_psum_27_50), .reg_activation(reg_activation_28_50), .reg_weight(reg_weight_28_50), .reg_partial_sum(reg_psum_28_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_51( .activation_in(reg_activation_28_50), .weight_in(reg_weight_27_51), .partial_sum_in(reg_psum_27_51), .reg_activation(reg_activation_28_51), .reg_weight(reg_weight_28_51), .reg_partial_sum(reg_psum_28_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_52( .activation_in(reg_activation_28_51), .weight_in(reg_weight_27_52), .partial_sum_in(reg_psum_27_52), .reg_activation(reg_activation_28_52), .reg_weight(reg_weight_28_52), .reg_partial_sum(reg_psum_28_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_53( .activation_in(reg_activation_28_52), .weight_in(reg_weight_27_53), .partial_sum_in(reg_psum_27_53), .reg_activation(reg_activation_28_53), .reg_weight(reg_weight_28_53), .reg_partial_sum(reg_psum_28_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_54( .activation_in(reg_activation_28_53), .weight_in(reg_weight_27_54), .partial_sum_in(reg_psum_27_54), .reg_activation(reg_activation_28_54), .reg_weight(reg_weight_28_54), .reg_partial_sum(reg_psum_28_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_55( .activation_in(reg_activation_28_54), .weight_in(reg_weight_27_55), .partial_sum_in(reg_psum_27_55), .reg_activation(reg_activation_28_55), .reg_weight(reg_weight_28_55), .reg_partial_sum(reg_psum_28_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_56( .activation_in(reg_activation_28_55), .weight_in(reg_weight_27_56), .partial_sum_in(reg_psum_27_56), .reg_activation(reg_activation_28_56), .reg_weight(reg_weight_28_56), .reg_partial_sum(reg_psum_28_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_57( .activation_in(reg_activation_28_56), .weight_in(reg_weight_27_57), .partial_sum_in(reg_psum_27_57), .reg_activation(reg_activation_28_57), .reg_weight(reg_weight_28_57), .reg_partial_sum(reg_psum_28_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_58( .activation_in(reg_activation_28_57), .weight_in(reg_weight_27_58), .partial_sum_in(reg_psum_27_58), .reg_activation(reg_activation_28_58), .reg_weight(reg_weight_28_58), .reg_partial_sum(reg_psum_28_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_59( .activation_in(reg_activation_28_58), .weight_in(reg_weight_27_59), .partial_sum_in(reg_psum_27_59), .reg_activation(reg_activation_28_59), .reg_weight(reg_weight_28_59), .reg_partial_sum(reg_psum_28_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_60( .activation_in(reg_activation_28_59), .weight_in(reg_weight_27_60), .partial_sum_in(reg_psum_27_60), .reg_activation(reg_activation_28_60), .reg_weight(reg_weight_28_60), .reg_partial_sum(reg_psum_28_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_61( .activation_in(reg_activation_28_60), .weight_in(reg_weight_27_61), .partial_sum_in(reg_psum_27_61), .reg_activation(reg_activation_28_61), .reg_weight(reg_weight_28_61), .reg_partial_sum(reg_psum_28_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_62( .activation_in(reg_activation_28_61), .weight_in(reg_weight_27_62), .partial_sum_in(reg_psum_27_62), .reg_activation(reg_activation_28_62), .reg_weight(reg_weight_28_62), .reg_partial_sum(reg_psum_28_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_63( .activation_in(reg_activation_28_62), .weight_in(reg_weight_27_63), .partial_sum_in(reg_psum_27_63), .reg_weight(reg_weight_28_63), .reg_partial_sum(reg_psum_28_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_0( .activation_in(in_activation_29), .weight_in(reg_weight_28_0), .partial_sum_in(reg_psum_28_0), .reg_activation(reg_activation_29_0), .reg_weight(reg_weight_29_0), .reg_partial_sum(reg_psum_29_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_1( .activation_in(reg_activation_29_0), .weight_in(reg_weight_28_1), .partial_sum_in(reg_psum_28_1), .reg_activation(reg_activation_29_1), .reg_weight(reg_weight_29_1), .reg_partial_sum(reg_psum_29_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_2( .activation_in(reg_activation_29_1), .weight_in(reg_weight_28_2), .partial_sum_in(reg_psum_28_2), .reg_activation(reg_activation_29_2), .reg_weight(reg_weight_29_2), .reg_partial_sum(reg_psum_29_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_3( .activation_in(reg_activation_29_2), .weight_in(reg_weight_28_3), .partial_sum_in(reg_psum_28_3), .reg_activation(reg_activation_29_3), .reg_weight(reg_weight_29_3), .reg_partial_sum(reg_psum_29_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_4( .activation_in(reg_activation_29_3), .weight_in(reg_weight_28_4), .partial_sum_in(reg_psum_28_4), .reg_activation(reg_activation_29_4), .reg_weight(reg_weight_29_4), .reg_partial_sum(reg_psum_29_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_5( .activation_in(reg_activation_29_4), .weight_in(reg_weight_28_5), .partial_sum_in(reg_psum_28_5), .reg_activation(reg_activation_29_5), .reg_weight(reg_weight_29_5), .reg_partial_sum(reg_psum_29_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_6( .activation_in(reg_activation_29_5), .weight_in(reg_weight_28_6), .partial_sum_in(reg_psum_28_6), .reg_activation(reg_activation_29_6), .reg_weight(reg_weight_29_6), .reg_partial_sum(reg_psum_29_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_7( .activation_in(reg_activation_29_6), .weight_in(reg_weight_28_7), .partial_sum_in(reg_psum_28_7), .reg_activation(reg_activation_29_7), .reg_weight(reg_weight_29_7), .reg_partial_sum(reg_psum_29_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_8( .activation_in(reg_activation_29_7), .weight_in(reg_weight_28_8), .partial_sum_in(reg_psum_28_8), .reg_activation(reg_activation_29_8), .reg_weight(reg_weight_29_8), .reg_partial_sum(reg_psum_29_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_9( .activation_in(reg_activation_29_8), .weight_in(reg_weight_28_9), .partial_sum_in(reg_psum_28_9), .reg_activation(reg_activation_29_9), .reg_weight(reg_weight_29_9), .reg_partial_sum(reg_psum_29_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_10( .activation_in(reg_activation_29_9), .weight_in(reg_weight_28_10), .partial_sum_in(reg_psum_28_10), .reg_activation(reg_activation_29_10), .reg_weight(reg_weight_29_10), .reg_partial_sum(reg_psum_29_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_11( .activation_in(reg_activation_29_10), .weight_in(reg_weight_28_11), .partial_sum_in(reg_psum_28_11), .reg_activation(reg_activation_29_11), .reg_weight(reg_weight_29_11), .reg_partial_sum(reg_psum_29_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_12( .activation_in(reg_activation_29_11), .weight_in(reg_weight_28_12), .partial_sum_in(reg_psum_28_12), .reg_activation(reg_activation_29_12), .reg_weight(reg_weight_29_12), .reg_partial_sum(reg_psum_29_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_13( .activation_in(reg_activation_29_12), .weight_in(reg_weight_28_13), .partial_sum_in(reg_psum_28_13), .reg_activation(reg_activation_29_13), .reg_weight(reg_weight_29_13), .reg_partial_sum(reg_psum_29_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_14( .activation_in(reg_activation_29_13), .weight_in(reg_weight_28_14), .partial_sum_in(reg_psum_28_14), .reg_activation(reg_activation_29_14), .reg_weight(reg_weight_29_14), .reg_partial_sum(reg_psum_29_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_15( .activation_in(reg_activation_29_14), .weight_in(reg_weight_28_15), .partial_sum_in(reg_psum_28_15), .reg_activation(reg_activation_29_15), .reg_weight(reg_weight_29_15), .reg_partial_sum(reg_psum_29_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_16( .activation_in(reg_activation_29_15), .weight_in(reg_weight_28_16), .partial_sum_in(reg_psum_28_16), .reg_activation(reg_activation_29_16), .reg_weight(reg_weight_29_16), .reg_partial_sum(reg_psum_29_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_17( .activation_in(reg_activation_29_16), .weight_in(reg_weight_28_17), .partial_sum_in(reg_psum_28_17), .reg_activation(reg_activation_29_17), .reg_weight(reg_weight_29_17), .reg_partial_sum(reg_psum_29_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_18( .activation_in(reg_activation_29_17), .weight_in(reg_weight_28_18), .partial_sum_in(reg_psum_28_18), .reg_activation(reg_activation_29_18), .reg_weight(reg_weight_29_18), .reg_partial_sum(reg_psum_29_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_19( .activation_in(reg_activation_29_18), .weight_in(reg_weight_28_19), .partial_sum_in(reg_psum_28_19), .reg_activation(reg_activation_29_19), .reg_weight(reg_weight_29_19), .reg_partial_sum(reg_psum_29_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_20( .activation_in(reg_activation_29_19), .weight_in(reg_weight_28_20), .partial_sum_in(reg_psum_28_20), .reg_activation(reg_activation_29_20), .reg_weight(reg_weight_29_20), .reg_partial_sum(reg_psum_29_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_21( .activation_in(reg_activation_29_20), .weight_in(reg_weight_28_21), .partial_sum_in(reg_psum_28_21), .reg_activation(reg_activation_29_21), .reg_weight(reg_weight_29_21), .reg_partial_sum(reg_psum_29_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_22( .activation_in(reg_activation_29_21), .weight_in(reg_weight_28_22), .partial_sum_in(reg_psum_28_22), .reg_activation(reg_activation_29_22), .reg_weight(reg_weight_29_22), .reg_partial_sum(reg_psum_29_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_23( .activation_in(reg_activation_29_22), .weight_in(reg_weight_28_23), .partial_sum_in(reg_psum_28_23), .reg_activation(reg_activation_29_23), .reg_weight(reg_weight_29_23), .reg_partial_sum(reg_psum_29_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_24( .activation_in(reg_activation_29_23), .weight_in(reg_weight_28_24), .partial_sum_in(reg_psum_28_24), .reg_activation(reg_activation_29_24), .reg_weight(reg_weight_29_24), .reg_partial_sum(reg_psum_29_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_25( .activation_in(reg_activation_29_24), .weight_in(reg_weight_28_25), .partial_sum_in(reg_psum_28_25), .reg_activation(reg_activation_29_25), .reg_weight(reg_weight_29_25), .reg_partial_sum(reg_psum_29_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_26( .activation_in(reg_activation_29_25), .weight_in(reg_weight_28_26), .partial_sum_in(reg_psum_28_26), .reg_activation(reg_activation_29_26), .reg_weight(reg_weight_29_26), .reg_partial_sum(reg_psum_29_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_27( .activation_in(reg_activation_29_26), .weight_in(reg_weight_28_27), .partial_sum_in(reg_psum_28_27), .reg_activation(reg_activation_29_27), .reg_weight(reg_weight_29_27), .reg_partial_sum(reg_psum_29_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_28( .activation_in(reg_activation_29_27), .weight_in(reg_weight_28_28), .partial_sum_in(reg_psum_28_28), .reg_activation(reg_activation_29_28), .reg_weight(reg_weight_29_28), .reg_partial_sum(reg_psum_29_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_29( .activation_in(reg_activation_29_28), .weight_in(reg_weight_28_29), .partial_sum_in(reg_psum_28_29), .reg_activation(reg_activation_29_29), .reg_weight(reg_weight_29_29), .reg_partial_sum(reg_psum_29_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_30( .activation_in(reg_activation_29_29), .weight_in(reg_weight_28_30), .partial_sum_in(reg_psum_28_30), .reg_activation(reg_activation_29_30), .reg_weight(reg_weight_29_30), .reg_partial_sum(reg_psum_29_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_31( .activation_in(reg_activation_29_30), .weight_in(reg_weight_28_31), .partial_sum_in(reg_psum_28_31), .reg_activation(reg_activation_29_31), .reg_weight(reg_weight_29_31), .reg_partial_sum(reg_psum_29_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_32( .activation_in(reg_activation_29_31), .weight_in(reg_weight_28_32), .partial_sum_in(reg_psum_28_32), .reg_activation(reg_activation_29_32), .reg_weight(reg_weight_29_32), .reg_partial_sum(reg_psum_29_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_33( .activation_in(reg_activation_29_32), .weight_in(reg_weight_28_33), .partial_sum_in(reg_psum_28_33), .reg_activation(reg_activation_29_33), .reg_weight(reg_weight_29_33), .reg_partial_sum(reg_psum_29_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_34( .activation_in(reg_activation_29_33), .weight_in(reg_weight_28_34), .partial_sum_in(reg_psum_28_34), .reg_activation(reg_activation_29_34), .reg_weight(reg_weight_29_34), .reg_partial_sum(reg_psum_29_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_35( .activation_in(reg_activation_29_34), .weight_in(reg_weight_28_35), .partial_sum_in(reg_psum_28_35), .reg_activation(reg_activation_29_35), .reg_weight(reg_weight_29_35), .reg_partial_sum(reg_psum_29_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_36( .activation_in(reg_activation_29_35), .weight_in(reg_weight_28_36), .partial_sum_in(reg_psum_28_36), .reg_activation(reg_activation_29_36), .reg_weight(reg_weight_29_36), .reg_partial_sum(reg_psum_29_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_37( .activation_in(reg_activation_29_36), .weight_in(reg_weight_28_37), .partial_sum_in(reg_psum_28_37), .reg_activation(reg_activation_29_37), .reg_weight(reg_weight_29_37), .reg_partial_sum(reg_psum_29_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_38( .activation_in(reg_activation_29_37), .weight_in(reg_weight_28_38), .partial_sum_in(reg_psum_28_38), .reg_activation(reg_activation_29_38), .reg_weight(reg_weight_29_38), .reg_partial_sum(reg_psum_29_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_39( .activation_in(reg_activation_29_38), .weight_in(reg_weight_28_39), .partial_sum_in(reg_psum_28_39), .reg_activation(reg_activation_29_39), .reg_weight(reg_weight_29_39), .reg_partial_sum(reg_psum_29_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_40( .activation_in(reg_activation_29_39), .weight_in(reg_weight_28_40), .partial_sum_in(reg_psum_28_40), .reg_activation(reg_activation_29_40), .reg_weight(reg_weight_29_40), .reg_partial_sum(reg_psum_29_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_41( .activation_in(reg_activation_29_40), .weight_in(reg_weight_28_41), .partial_sum_in(reg_psum_28_41), .reg_activation(reg_activation_29_41), .reg_weight(reg_weight_29_41), .reg_partial_sum(reg_psum_29_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_42( .activation_in(reg_activation_29_41), .weight_in(reg_weight_28_42), .partial_sum_in(reg_psum_28_42), .reg_activation(reg_activation_29_42), .reg_weight(reg_weight_29_42), .reg_partial_sum(reg_psum_29_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_43( .activation_in(reg_activation_29_42), .weight_in(reg_weight_28_43), .partial_sum_in(reg_psum_28_43), .reg_activation(reg_activation_29_43), .reg_weight(reg_weight_29_43), .reg_partial_sum(reg_psum_29_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_44( .activation_in(reg_activation_29_43), .weight_in(reg_weight_28_44), .partial_sum_in(reg_psum_28_44), .reg_activation(reg_activation_29_44), .reg_weight(reg_weight_29_44), .reg_partial_sum(reg_psum_29_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_45( .activation_in(reg_activation_29_44), .weight_in(reg_weight_28_45), .partial_sum_in(reg_psum_28_45), .reg_activation(reg_activation_29_45), .reg_weight(reg_weight_29_45), .reg_partial_sum(reg_psum_29_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_46( .activation_in(reg_activation_29_45), .weight_in(reg_weight_28_46), .partial_sum_in(reg_psum_28_46), .reg_activation(reg_activation_29_46), .reg_weight(reg_weight_29_46), .reg_partial_sum(reg_psum_29_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_47( .activation_in(reg_activation_29_46), .weight_in(reg_weight_28_47), .partial_sum_in(reg_psum_28_47), .reg_activation(reg_activation_29_47), .reg_weight(reg_weight_29_47), .reg_partial_sum(reg_psum_29_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_48( .activation_in(reg_activation_29_47), .weight_in(reg_weight_28_48), .partial_sum_in(reg_psum_28_48), .reg_activation(reg_activation_29_48), .reg_weight(reg_weight_29_48), .reg_partial_sum(reg_psum_29_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_49( .activation_in(reg_activation_29_48), .weight_in(reg_weight_28_49), .partial_sum_in(reg_psum_28_49), .reg_activation(reg_activation_29_49), .reg_weight(reg_weight_29_49), .reg_partial_sum(reg_psum_29_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_50( .activation_in(reg_activation_29_49), .weight_in(reg_weight_28_50), .partial_sum_in(reg_psum_28_50), .reg_activation(reg_activation_29_50), .reg_weight(reg_weight_29_50), .reg_partial_sum(reg_psum_29_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_51( .activation_in(reg_activation_29_50), .weight_in(reg_weight_28_51), .partial_sum_in(reg_psum_28_51), .reg_activation(reg_activation_29_51), .reg_weight(reg_weight_29_51), .reg_partial_sum(reg_psum_29_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_52( .activation_in(reg_activation_29_51), .weight_in(reg_weight_28_52), .partial_sum_in(reg_psum_28_52), .reg_activation(reg_activation_29_52), .reg_weight(reg_weight_29_52), .reg_partial_sum(reg_psum_29_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_53( .activation_in(reg_activation_29_52), .weight_in(reg_weight_28_53), .partial_sum_in(reg_psum_28_53), .reg_activation(reg_activation_29_53), .reg_weight(reg_weight_29_53), .reg_partial_sum(reg_psum_29_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_54( .activation_in(reg_activation_29_53), .weight_in(reg_weight_28_54), .partial_sum_in(reg_psum_28_54), .reg_activation(reg_activation_29_54), .reg_weight(reg_weight_29_54), .reg_partial_sum(reg_psum_29_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_55( .activation_in(reg_activation_29_54), .weight_in(reg_weight_28_55), .partial_sum_in(reg_psum_28_55), .reg_activation(reg_activation_29_55), .reg_weight(reg_weight_29_55), .reg_partial_sum(reg_psum_29_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_56( .activation_in(reg_activation_29_55), .weight_in(reg_weight_28_56), .partial_sum_in(reg_psum_28_56), .reg_activation(reg_activation_29_56), .reg_weight(reg_weight_29_56), .reg_partial_sum(reg_psum_29_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_57( .activation_in(reg_activation_29_56), .weight_in(reg_weight_28_57), .partial_sum_in(reg_psum_28_57), .reg_activation(reg_activation_29_57), .reg_weight(reg_weight_29_57), .reg_partial_sum(reg_psum_29_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_58( .activation_in(reg_activation_29_57), .weight_in(reg_weight_28_58), .partial_sum_in(reg_psum_28_58), .reg_activation(reg_activation_29_58), .reg_weight(reg_weight_29_58), .reg_partial_sum(reg_psum_29_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_59( .activation_in(reg_activation_29_58), .weight_in(reg_weight_28_59), .partial_sum_in(reg_psum_28_59), .reg_activation(reg_activation_29_59), .reg_weight(reg_weight_29_59), .reg_partial_sum(reg_psum_29_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_60( .activation_in(reg_activation_29_59), .weight_in(reg_weight_28_60), .partial_sum_in(reg_psum_28_60), .reg_activation(reg_activation_29_60), .reg_weight(reg_weight_29_60), .reg_partial_sum(reg_psum_29_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_61( .activation_in(reg_activation_29_60), .weight_in(reg_weight_28_61), .partial_sum_in(reg_psum_28_61), .reg_activation(reg_activation_29_61), .reg_weight(reg_weight_29_61), .reg_partial_sum(reg_psum_29_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_62( .activation_in(reg_activation_29_61), .weight_in(reg_weight_28_62), .partial_sum_in(reg_psum_28_62), .reg_activation(reg_activation_29_62), .reg_weight(reg_weight_29_62), .reg_partial_sum(reg_psum_29_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_63( .activation_in(reg_activation_29_62), .weight_in(reg_weight_28_63), .partial_sum_in(reg_psum_28_63), .reg_weight(reg_weight_29_63), .reg_partial_sum(reg_psum_29_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_0( .activation_in(in_activation_30), .weight_in(reg_weight_29_0), .partial_sum_in(reg_psum_29_0), .reg_activation(reg_activation_30_0), .reg_weight(reg_weight_30_0), .reg_partial_sum(reg_psum_30_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_1( .activation_in(reg_activation_30_0), .weight_in(reg_weight_29_1), .partial_sum_in(reg_psum_29_1), .reg_activation(reg_activation_30_1), .reg_weight(reg_weight_30_1), .reg_partial_sum(reg_psum_30_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_2( .activation_in(reg_activation_30_1), .weight_in(reg_weight_29_2), .partial_sum_in(reg_psum_29_2), .reg_activation(reg_activation_30_2), .reg_weight(reg_weight_30_2), .reg_partial_sum(reg_psum_30_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_3( .activation_in(reg_activation_30_2), .weight_in(reg_weight_29_3), .partial_sum_in(reg_psum_29_3), .reg_activation(reg_activation_30_3), .reg_weight(reg_weight_30_3), .reg_partial_sum(reg_psum_30_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_4( .activation_in(reg_activation_30_3), .weight_in(reg_weight_29_4), .partial_sum_in(reg_psum_29_4), .reg_activation(reg_activation_30_4), .reg_weight(reg_weight_30_4), .reg_partial_sum(reg_psum_30_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_5( .activation_in(reg_activation_30_4), .weight_in(reg_weight_29_5), .partial_sum_in(reg_psum_29_5), .reg_activation(reg_activation_30_5), .reg_weight(reg_weight_30_5), .reg_partial_sum(reg_psum_30_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_6( .activation_in(reg_activation_30_5), .weight_in(reg_weight_29_6), .partial_sum_in(reg_psum_29_6), .reg_activation(reg_activation_30_6), .reg_weight(reg_weight_30_6), .reg_partial_sum(reg_psum_30_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_7( .activation_in(reg_activation_30_6), .weight_in(reg_weight_29_7), .partial_sum_in(reg_psum_29_7), .reg_activation(reg_activation_30_7), .reg_weight(reg_weight_30_7), .reg_partial_sum(reg_psum_30_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_8( .activation_in(reg_activation_30_7), .weight_in(reg_weight_29_8), .partial_sum_in(reg_psum_29_8), .reg_activation(reg_activation_30_8), .reg_weight(reg_weight_30_8), .reg_partial_sum(reg_psum_30_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_9( .activation_in(reg_activation_30_8), .weight_in(reg_weight_29_9), .partial_sum_in(reg_psum_29_9), .reg_activation(reg_activation_30_9), .reg_weight(reg_weight_30_9), .reg_partial_sum(reg_psum_30_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_10( .activation_in(reg_activation_30_9), .weight_in(reg_weight_29_10), .partial_sum_in(reg_psum_29_10), .reg_activation(reg_activation_30_10), .reg_weight(reg_weight_30_10), .reg_partial_sum(reg_psum_30_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_11( .activation_in(reg_activation_30_10), .weight_in(reg_weight_29_11), .partial_sum_in(reg_psum_29_11), .reg_activation(reg_activation_30_11), .reg_weight(reg_weight_30_11), .reg_partial_sum(reg_psum_30_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_12( .activation_in(reg_activation_30_11), .weight_in(reg_weight_29_12), .partial_sum_in(reg_psum_29_12), .reg_activation(reg_activation_30_12), .reg_weight(reg_weight_30_12), .reg_partial_sum(reg_psum_30_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_13( .activation_in(reg_activation_30_12), .weight_in(reg_weight_29_13), .partial_sum_in(reg_psum_29_13), .reg_activation(reg_activation_30_13), .reg_weight(reg_weight_30_13), .reg_partial_sum(reg_psum_30_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_14( .activation_in(reg_activation_30_13), .weight_in(reg_weight_29_14), .partial_sum_in(reg_psum_29_14), .reg_activation(reg_activation_30_14), .reg_weight(reg_weight_30_14), .reg_partial_sum(reg_psum_30_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_15( .activation_in(reg_activation_30_14), .weight_in(reg_weight_29_15), .partial_sum_in(reg_psum_29_15), .reg_activation(reg_activation_30_15), .reg_weight(reg_weight_30_15), .reg_partial_sum(reg_psum_30_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_16( .activation_in(reg_activation_30_15), .weight_in(reg_weight_29_16), .partial_sum_in(reg_psum_29_16), .reg_activation(reg_activation_30_16), .reg_weight(reg_weight_30_16), .reg_partial_sum(reg_psum_30_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_17( .activation_in(reg_activation_30_16), .weight_in(reg_weight_29_17), .partial_sum_in(reg_psum_29_17), .reg_activation(reg_activation_30_17), .reg_weight(reg_weight_30_17), .reg_partial_sum(reg_psum_30_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_18( .activation_in(reg_activation_30_17), .weight_in(reg_weight_29_18), .partial_sum_in(reg_psum_29_18), .reg_activation(reg_activation_30_18), .reg_weight(reg_weight_30_18), .reg_partial_sum(reg_psum_30_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_19( .activation_in(reg_activation_30_18), .weight_in(reg_weight_29_19), .partial_sum_in(reg_psum_29_19), .reg_activation(reg_activation_30_19), .reg_weight(reg_weight_30_19), .reg_partial_sum(reg_psum_30_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_20( .activation_in(reg_activation_30_19), .weight_in(reg_weight_29_20), .partial_sum_in(reg_psum_29_20), .reg_activation(reg_activation_30_20), .reg_weight(reg_weight_30_20), .reg_partial_sum(reg_psum_30_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_21( .activation_in(reg_activation_30_20), .weight_in(reg_weight_29_21), .partial_sum_in(reg_psum_29_21), .reg_activation(reg_activation_30_21), .reg_weight(reg_weight_30_21), .reg_partial_sum(reg_psum_30_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_22( .activation_in(reg_activation_30_21), .weight_in(reg_weight_29_22), .partial_sum_in(reg_psum_29_22), .reg_activation(reg_activation_30_22), .reg_weight(reg_weight_30_22), .reg_partial_sum(reg_psum_30_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_23( .activation_in(reg_activation_30_22), .weight_in(reg_weight_29_23), .partial_sum_in(reg_psum_29_23), .reg_activation(reg_activation_30_23), .reg_weight(reg_weight_30_23), .reg_partial_sum(reg_psum_30_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_24( .activation_in(reg_activation_30_23), .weight_in(reg_weight_29_24), .partial_sum_in(reg_psum_29_24), .reg_activation(reg_activation_30_24), .reg_weight(reg_weight_30_24), .reg_partial_sum(reg_psum_30_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_25( .activation_in(reg_activation_30_24), .weight_in(reg_weight_29_25), .partial_sum_in(reg_psum_29_25), .reg_activation(reg_activation_30_25), .reg_weight(reg_weight_30_25), .reg_partial_sum(reg_psum_30_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_26( .activation_in(reg_activation_30_25), .weight_in(reg_weight_29_26), .partial_sum_in(reg_psum_29_26), .reg_activation(reg_activation_30_26), .reg_weight(reg_weight_30_26), .reg_partial_sum(reg_psum_30_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_27( .activation_in(reg_activation_30_26), .weight_in(reg_weight_29_27), .partial_sum_in(reg_psum_29_27), .reg_activation(reg_activation_30_27), .reg_weight(reg_weight_30_27), .reg_partial_sum(reg_psum_30_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_28( .activation_in(reg_activation_30_27), .weight_in(reg_weight_29_28), .partial_sum_in(reg_psum_29_28), .reg_activation(reg_activation_30_28), .reg_weight(reg_weight_30_28), .reg_partial_sum(reg_psum_30_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_29( .activation_in(reg_activation_30_28), .weight_in(reg_weight_29_29), .partial_sum_in(reg_psum_29_29), .reg_activation(reg_activation_30_29), .reg_weight(reg_weight_30_29), .reg_partial_sum(reg_psum_30_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_30( .activation_in(reg_activation_30_29), .weight_in(reg_weight_29_30), .partial_sum_in(reg_psum_29_30), .reg_activation(reg_activation_30_30), .reg_weight(reg_weight_30_30), .reg_partial_sum(reg_psum_30_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_31( .activation_in(reg_activation_30_30), .weight_in(reg_weight_29_31), .partial_sum_in(reg_psum_29_31), .reg_activation(reg_activation_30_31), .reg_weight(reg_weight_30_31), .reg_partial_sum(reg_psum_30_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_32( .activation_in(reg_activation_30_31), .weight_in(reg_weight_29_32), .partial_sum_in(reg_psum_29_32), .reg_activation(reg_activation_30_32), .reg_weight(reg_weight_30_32), .reg_partial_sum(reg_psum_30_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_33( .activation_in(reg_activation_30_32), .weight_in(reg_weight_29_33), .partial_sum_in(reg_psum_29_33), .reg_activation(reg_activation_30_33), .reg_weight(reg_weight_30_33), .reg_partial_sum(reg_psum_30_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_34( .activation_in(reg_activation_30_33), .weight_in(reg_weight_29_34), .partial_sum_in(reg_psum_29_34), .reg_activation(reg_activation_30_34), .reg_weight(reg_weight_30_34), .reg_partial_sum(reg_psum_30_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_35( .activation_in(reg_activation_30_34), .weight_in(reg_weight_29_35), .partial_sum_in(reg_psum_29_35), .reg_activation(reg_activation_30_35), .reg_weight(reg_weight_30_35), .reg_partial_sum(reg_psum_30_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_36( .activation_in(reg_activation_30_35), .weight_in(reg_weight_29_36), .partial_sum_in(reg_psum_29_36), .reg_activation(reg_activation_30_36), .reg_weight(reg_weight_30_36), .reg_partial_sum(reg_psum_30_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_37( .activation_in(reg_activation_30_36), .weight_in(reg_weight_29_37), .partial_sum_in(reg_psum_29_37), .reg_activation(reg_activation_30_37), .reg_weight(reg_weight_30_37), .reg_partial_sum(reg_psum_30_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_38( .activation_in(reg_activation_30_37), .weight_in(reg_weight_29_38), .partial_sum_in(reg_psum_29_38), .reg_activation(reg_activation_30_38), .reg_weight(reg_weight_30_38), .reg_partial_sum(reg_psum_30_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_39( .activation_in(reg_activation_30_38), .weight_in(reg_weight_29_39), .partial_sum_in(reg_psum_29_39), .reg_activation(reg_activation_30_39), .reg_weight(reg_weight_30_39), .reg_partial_sum(reg_psum_30_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_40( .activation_in(reg_activation_30_39), .weight_in(reg_weight_29_40), .partial_sum_in(reg_psum_29_40), .reg_activation(reg_activation_30_40), .reg_weight(reg_weight_30_40), .reg_partial_sum(reg_psum_30_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_41( .activation_in(reg_activation_30_40), .weight_in(reg_weight_29_41), .partial_sum_in(reg_psum_29_41), .reg_activation(reg_activation_30_41), .reg_weight(reg_weight_30_41), .reg_partial_sum(reg_psum_30_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_42( .activation_in(reg_activation_30_41), .weight_in(reg_weight_29_42), .partial_sum_in(reg_psum_29_42), .reg_activation(reg_activation_30_42), .reg_weight(reg_weight_30_42), .reg_partial_sum(reg_psum_30_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_43( .activation_in(reg_activation_30_42), .weight_in(reg_weight_29_43), .partial_sum_in(reg_psum_29_43), .reg_activation(reg_activation_30_43), .reg_weight(reg_weight_30_43), .reg_partial_sum(reg_psum_30_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_44( .activation_in(reg_activation_30_43), .weight_in(reg_weight_29_44), .partial_sum_in(reg_psum_29_44), .reg_activation(reg_activation_30_44), .reg_weight(reg_weight_30_44), .reg_partial_sum(reg_psum_30_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_45( .activation_in(reg_activation_30_44), .weight_in(reg_weight_29_45), .partial_sum_in(reg_psum_29_45), .reg_activation(reg_activation_30_45), .reg_weight(reg_weight_30_45), .reg_partial_sum(reg_psum_30_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_46( .activation_in(reg_activation_30_45), .weight_in(reg_weight_29_46), .partial_sum_in(reg_psum_29_46), .reg_activation(reg_activation_30_46), .reg_weight(reg_weight_30_46), .reg_partial_sum(reg_psum_30_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_47( .activation_in(reg_activation_30_46), .weight_in(reg_weight_29_47), .partial_sum_in(reg_psum_29_47), .reg_activation(reg_activation_30_47), .reg_weight(reg_weight_30_47), .reg_partial_sum(reg_psum_30_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_48( .activation_in(reg_activation_30_47), .weight_in(reg_weight_29_48), .partial_sum_in(reg_psum_29_48), .reg_activation(reg_activation_30_48), .reg_weight(reg_weight_30_48), .reg_partial_sum(reg_psum_30_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_49( .activation_in(reg_activation_30_48), .weight_in(reg_weight_29_49), .partial_sum_in(reg_psum_29_49), .reg_activation(reg_activation_30_49), .reg_weight(reg_weight_30_49), .reg_partial_sum(reg_psum_30_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_50( .activation_in(reg_activation_30_49), .weight_in(reg_weight_29_50), .partial_sum_in(reg_psum_29_50), .reg_activation(reg_activation_30_50), .reg_weight(reg_weight_30_50), .reg_partial_sum(reg_psum_30_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_51( .activation_in(reg_activation_30_50), .weight_in(reg_weight_29_51), .partial_sum_in(reg_psum_29_51), .reg_activation(reg_activation_30_51), .reg_weight(reg_weight_30_51), .reg_partial_sum(reg_psum_30_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_52( .activation_in(reg_activation_30_51), .weight_in(reg_weight_29_52), .partial_sum_in(reg_psum_29_52), .reg_activation(reg_activation_30_52), .reg_weight(reg_weight_30_52), .reg_partial_sum(reg_psum_30_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_53( .activation_in(reg_activation_30_52), .weight_in(reg_weight_29_53), .partial_sum_in(reg_psum_29_53), .reg_activation(reg_activation_30_53), .reg_weight(reg_weight_30_53), .reg_partial_sum(reg_psum_30_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_54( .activation_in(reg_activation_30_53), .weight_in(reg_weight_29_54), .partial_sum_in(reg_psum_29_54), .reg_activation(reg_activation_30_54), .reg_weight(reg_weight_30_54), .reg_partial_sum(reg_psum_30_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_55( .activation_in(reg_activation_30_54), .weight_in(reg_weight_29_55), .partial_sum_in(reg_psum_29_55), .reg_activation(reg_activation_30_55), .reg_weight(reg_weight_30_55), .reg_partial_sum(reg_psum_30_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_56( .activation_in(reg_activation_30_55), .weight_in(reg_weight_29_56), .partial_sum_in(reg_psum_29_56), .reg_activation(reg_activation_30_56), .reg_weight(reg_weight_30_56), .reg_partial_sum(reg_psum_30_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_57( .activation_in(reg_activation_30_56), .weight_in(reg_weight_29_57), .partial_sum_in(reg_psum_29_57), .reg_activation(reg_activation_30_57), .reg_weight(reg_weight_30_57), .reg_partial_sum(reg_psum_30_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_58( .activation_in(reg_activation_30_57), .weight_in(reg_weight_29_58), .partial_sum_in(reg_psum_29_58), .reg_activation(reg_activation_30_58), .reg_weight(reg_weight_30_58), .reg_partial_sum(reg_psum_30_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_59( .activation_in(reg_activation_30_58), .weight_in(reg_weight_29_59), .partial_sum_in(reg_psum_29_59), .reg_activation(reg_activation_30_59), .reg_weight(reg_weight_30_59), .reg_partial_sum(reg_psum_30_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_60( .activation_in(reg_activation_30_59), .weight_in(reg_weight_29_60), .partial_sum_in(reg_psum_29_60), .reg_activation(reg_activation_30_60), .reg_weight(reg_weight_30_60), .reg_partial_sum(reg_psum_30_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_61( .activation_in(reg_activation_30_60), .weight_in(reg_weight_29_61), .partial_sum_in(reg_psum_29_61), .reg_activation(reg_activation_30_61), .reg_weight(reg_weight_30_61), .reg_partial_sum(reg_psum_30_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_62( .activation_in(reg_activation_30_61), .weight_in(reg_weight_29_62), .partial_sum_in(reg_psum_29_62), .reg_activation(reg_activation_30_62), .reg_weight(reg_weight_30_62), .reg_partial_sum(reg_psum_30_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_63( .activation_in(reg_activation_30_62), .weight_in(reg_weight_29_63), .partial_sum_in(reg_psum_29_63), .reg_weight(reg_weight_30_63), .reg_partial_sum(reg_psum_30_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_0( .activation_in(in_activation_31), .weight_in(reg_weight_30_0), .partial_sum_in(reg_psum_30_0), .reg_activation(reg_activation_31_0), .reg_weight(reg_weight_31_0), .reg_partial_sum(reg_psum_31_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_1( .activation_in(reg_activation_31_0), .weight_in(reg_weight_30_1), .partial_sum_in(reg_psum_30_1), .reg_activation(reg_activation_31_1), .reg_weight(reg_weight_31_1), .reg_partial_sum(reg_psum_31_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_2( .activation_in(reg_activation_31_1), .weight_in(reg_weight_30_2), .partial_sum_in(reg_psum_30_2), .reg_activation(reg_activation_31_2), .reg_weight(reg_weight_31_2), .reg_partial_sum(reg_psum_31_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_3( .activation_in(reg_activation_31_2), .weight_in(reg_weight_30_3), .partial_sum_in(reg_psum_30_3), .reg_activation(reg_activation_31_3), .reg_weight(reg_weight_31_3), .reg_partial_sum(reg_psum_31_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_4( .activation_in(reg_activation_31_3), .weight_in(reg_weight_30_4), .partial_sum_in(reg_psum_30_4), .reg_activation(reg_activation_31_4), .reg_weight(reg_weight_31_4), .reg_partial_sum(reg_psum_31_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_5( .activation_in(reg_activation_31_4), .weight_in(reg_weight_30_5), .partial_sum_in(reg_psum_30_5), .reg_activation(reg_activation_31_5), .reg_weight(reg_weight_31_5), .reg_partial_sum(reg_psum_31_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_6( .activation_in(reg_activation_31_5), .weight_in(reg_weight_30_6), .partial_sum_in(reg_psum_30_6), .reg_activation(reg_activation_31_6), .reg_weight(reg_weight_31_6), .reg_partial_sum(reg_psum_31_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_7( .activation_in(reg_activation_31_6), .weight_in(reg_weight_30_7), .partial_sum_in(reg_psum_30_7), .reg_activation(reg_activation_31_7), .reg_weight(reg_weight_31_7), .reg_partial_sum(reg_psum_31_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_8( .activation_in(reg_activation_31_7), .weight_in(reg_weight_30_8), .partial_sum_in(reg_psum_30_8), .reg_activation(reg_activation_31_8), .reg_weight(reg_weight_31_8), .reg_partial_sum(reg_psum_31_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_9( .activation_in(reg_activation_31_8), .weight_in(reg_weight_30_9), .partial_sum_in(reg_psum_30_9), .reg_activation(reg_activation_31_9), .reg_weight(reg_weight_31_9), .reg_partial_sum(reg_psum_31_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_10( .activation_in(reg_activation_31_9), .weight_in(reg_weight_30_10), .partial_sum_in(reg_psum_30_10), .reg_activation(reg_activation_31_10), .reg_weight(reg_weight_31_10), .reg_partial_sum(reg_psum_31_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_11( .activation_in(reg_activation_31_10), .weight_in(reg_weight_30_11), .partial_sum_in(reg_psum_30_11), .reg_activation(reg_activation_31_11), .reg_weight(reg_weight_31_11), .reg_partial_sum(reg_psum_31_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_12( .activation_in(reg_activation_31_11), .weight_in(reg_weight_30_12), .partial_sum_in(reg_psum_30_12), .reg_activation(reg_activation_31_12), .reg_weight(reg_weight_31_12), .reg_partial_sum(reg_psum_31_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_13( .activation_in(reg_activation_31_12), .weight_in(reg_weight_30_13), .partial_sum_in(reg_psum_30_13), .reg_activation(reg_activation_31_13), .reg_weight(reg_weight_31_13), .reg_partial_sum(reg_psum_31_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_14( .activation_in(reg_activation_31_13), .weight_in(reg_weight_30_14), .partial_sum_in(reg_psum_30_14), .reg_activation(reg_activation_31_14), .reg_weight(reg_weight_31_14), .reg_partial_sum(reg_psum_31_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_15( .activation_in(reg_activation_31_14), .weight_in(reg_weight_30_15), .partial_sum_in(reg_psum_30_15), .reg_activation(reg_activation_31_15), .reg_weight(reg_weight_31_15), .reg_partial_sum(reg_psum_31_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_16( .activation_in(reg_activation_31_15), .weight_in(reg_weight_30_16), .partial_sum_in(reg_psum_30_16), .reg_activation(reg_activation_31_16), .reg_weight(reg_weight_31_16), .reg_partial_sum(reg_psum_31_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_17( .activation_in(reg_activation_31_16), .weight_in(reg_weight_30_17), .partial_sum_in(reg_psum_30_17), .reg_activation(reg_activation_31_17), .reg_weight(reg_weight_31_17), .reg_partial_sum(reg_psum_31_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_18( .activation_in(reg_activation_31_17), .weight_in(reg_weight_30_18), .partial_sum_in(reg_psum_30_18), .reg_activation(reg_activation_31_18), .reg_weight(reg_weight_31_18), .reg_partial_sum(reg_psum_31_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_19( .activation_in(reg_activation_31_18), .weight_in(reg_weight_30_19), .partial_sum_in(reg_psum_30_19), .reg_activation(reg_activation_31_19), .reg_weight(reg_weight_31_19), .reg_partial_sum(reg_psum_31_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_20( .activation_in(reg_activation_31_19), .weight_in(reg_weight_30_20), .partial_sum_in(reg_psum_30_20), .reg_activation(reg_activation_31_20), .reg_weight(reg_weight_31_20), .reg_partial_sum(reg_psum_31_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_21( .activation_in(reg_activation_31_20), .weight_in(reg_weight_30_21), .partial_sum_in(reg_psum_30_21), .reg_activation(reg_activation_31_21), .reg_weight(reg_weight_31_21), .reg_partial_sum(reg_psum_31_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_22( .activation_in(reg_activation_31_21), .weight_in(reg_weight_30_22), .partial_sum_in(reg_psum_30_22), .reg_activation(reg_activation_31_22), .reg_weight(reg_weight_31_22), .reg_partial_sum(reg_psum_31_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_23( .activation_in(reg_activation_31_22), .weight_in(reg_weight_30_23), .partial_sum_in(reg_psum_30_23), .reg_activation(reg_activation_31_23), .reg_weight(reg_weight_31_23), .reg_partial_sum(reg_psum_31_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_24( .activation_in(reg_activation_31_23), .weight_in(reg_weight_30_24), .partial_sum_in(reg_psum_30_24), .reg_activation(reg_activation_31_24), .reg_weight(reg_weight_31_24), .reg_partial_sum(reg_psum_31_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_25( .activation_in(reg_activation_31_24), .weight_in(reg_weight_30_25), .partial_sum_in(reg_psum_30_25), .reg_activation(reg_activation_31_25), .reg_weight(reg_weight_31_25), .reg_partial_sum(reg_psum_31_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_26( .activation_in(reg_activation_31_25), .weight_in(reg_weight_30_26), .partial_sum_in(reg_psum_30_26), .reg_activation(reg_activation_31_26), .reg_weight(reg_weight_31_26), .reg_partial_sum(reg_psum_31_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_27( .activation_in(reg_activation_31_26), .weight_in(reg_weight_30_27), .partial_sum_in(reg_psum_30_27), .reg_activation(reg_activation_31_27), .reg_weight(reg_weight_31_27), .reg_partial_sum(reg_psum_31_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_28( .activation_in(reg_activation_31_27), .weight_in(reg_weight_30_28), .partial_sum_in(reg_psum_30_28), .reg_activation(reg_activation_31_28), .reg_weight(reg_weight_31_28), .reg_partial_sum(reg_psum_31_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_29( .activation_in(reg_activation_31_28), .weight_in(reg_weight_30_29), .partial_sum_in(reg_psum_30_29), .reg_activation(reg_activation_31_29), .reg_weight(reg_weight_31_29), .reg_partial_sum(reg_psum_31_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_30( .activation_in(reg_activation_31_29), .weight_in(reg_weight_30_30), .partial_sum_in(reg_psum_30_30), .reg_activation(reg_activation_31_30), .reg_weight(reg_weight_31_30), .reg_partial_sum(reg_psum_31_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_31( .activation_in(reg_activation_31_30), .weight_in(reg_weight_30_31), .partial_sum_in(reg_psum_30_31), .reg_activation(reg_activation_31_31), .reg_weight(reg_weight_31_31), .reg_partial_sum(reg_psum_31_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_32( .activation_in(reg_activation_31_31), .weight_in(reg_weight_30_32), .partial_sum_in(reg_psum_30_32), .reg_activation(reg_activation_31_32), .reg_weight(reg_weight_31_32), .reg_partial_sum(reg_psum_31_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_33( .activation_in(reg_activation_31_32), .weight_in(reg_weight_30_33), .partial_sum_in(reg_psum_30_33), .reg_activation(reg_activation_31_33), .reg_weight(reg_weight_31_33), .reg_partial_sum(reg_psum_31_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_34( .activation_in(reg_activation_31_33), .weight_in(reg_weight_30_34), .partial_sum_in(reg_psum_30_34), .reg_activation(reg_activation_31_34), .reg_weight(reg_weight_31_34), .reg_partial_sum(reg_psum_31_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_35( .activation_in(reg_activation_31_34), .weight_in(reg_weight_30_35), .partial_sum_in(reg_psum_30_35), .reg_activation(reg_activation_31_35), .reg_weight(reg_weight_31_35), .reg_partial_sum(reg_psum_31_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_36( .activation_in(reg_activation_31_35), .weight_in(reg_weight_30_36), .partial_sum_in(reg_psum_30_36), .reg_activation(reg_activation_31_36), .reg_weight(reg_weight_31_36), .reg_partial_sum(reg_psum_31_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_37( .activation_in(reg_activation_31_36), .weight_in(reg_weight_30_37), .partial_sum_in(reg_psum_30_37), .reg_activation(reg_activation_31_37), .reg_weight(reg_weight_31_37), .reg_partial_sum(reg_psum_31_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_38( .activation_in(reg_activation_31_37), .weight_in(reg_weight_30_38), .partial_sum_in(reg_psum_30_38), .reg_activation(reg_activation_31_38), .reg_weight(reg_weight_31_38), .reg_partial_sum(reg_psum_31_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_39( .activation_in(reg_activation_31_38), .weight_in(reg_weight_30_39), .partial_sum_in(reg_psum_30_39), .reg_activation(reg_activation_31_39), .reg_weight(reg_weight_31_39), .reg_partial_sum(reg_psum_31_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_40( .activation_in(reg_activation_31_39), .weight_in(reg_weight_30_40), .partial_sum_in(reg_psum_30_40), .reg_activation(reg_activation_31_40), .reg_weight(reg_weight_31_40), .reg_partial_sum(reg_psum_31_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_41( .activation_in(reg_activation_31_40), .weight_in(reg_weight_30_41), .partial_sum_in(reg_psum_30_41), .reg_activation(reg_activation_31_41), .reg_weight(reg_weight_31_41), .reg_partial_sum(reg_psum_31_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_42( .activation_in(reg_activation_31_41), .weight_in(reg_weight_30_42), .partial_sum_in(reg_psum_30_42), .reg_activation(reg_activation_31_42), .reg_weight(reg_weight_31_42), .reg_partial_sum(reg_psum_31_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_43( .activation_in(reg_activation_31_42), .weight_in(reg_weight_30_43), .partial_sum_in(reg_psum_30_43), .reg_activation(reg_activation_31_43), .reg_weight(reg_weight_31_43), .reg_partial_sum(reg_psum_31_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_44( .activation_in(reg_activation_31_43), .weight_in(reg_weight_30_44), .partial_sum_in(reg_psum_30_44), .reg_activation(reg_activation_31_44), .reg_weight(reg_weight_31_44), .reg_partial_sum(reg_psum_31_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_45( .activation_in(reg_activation_31_44), .weight_in(reg_weight_30_45), .partial_sum_in(reg_psum_30_45), .reg_activation(reg_activation_31_45), .reg_weight(reg_weight_31_45), .reg_partial_sum(reg_psum_31_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_46( .activation_in(reg_activation_31_45), .weight_in(reg_weight_30_46), .partial_sum_in(reg_psum_30_46), .reg_activation(reg_activation_31_46), .reg_weight(reg_weight_31_46), .reg_partial_sum(reg_psum_31_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_47( .activation_in(reg_activation_31_46), .weight_in(reg_weight_30_47), .partial_sum_in(reg_psum_30_47), .reg_activation(reg_activation_31_47), .reg_weight(reg_weight_31_47), .reg_partial_sum(reg_psum_31_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_48( .activation_in(reg_activation_31_47), .weight_in(reg_weight_30_48), .partial_sum_in(reg_psum_30_48), .reg_activation(reg_activation_31_48), .reg_weight(reg_weight_31_48), .reg_partial_sum(reg_psum_31_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_49( .activation_in(reg_activation_31_48), .weight_in(reg_weight_30_49), .partial_sum_in(reg_psum_30_49), .reg_activation(reg_activation_31_49), .reg_weight(reg_weight_31_49), .reg_partial_sum(reg_psum_31_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_50( .activation_in(reg_activation_31_49), .weight_in(reg_weight_30_50), .partial_sum_in(reg_psum_30_50), .reg_activation(reg_activation_31_50), .reg_weight(reg_weight_31_50), .reg_partial_sum(reg_psum_31_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_51( .activation_in(reg_activation_31_50), .weight_in(reg_weight_30_51), .partial_sum_in(reg_psum_30_51), .reg_activation(reg_activation_31_51), .reg_weight(reg_weight_31_51), .reg_partial_sum(reg_psum_31_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_52( .activation_in(reg_activation_31_51), .weight_in(reg_weight_30_52), .partial_sum_in(reg_psum_30_52), .reg_activation(reg_activation_31_52), .reg_weight(reg_weight_31_52), .reg_partial_sum(reg_psum_31_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_53( .activation_in(reg_activation_31_52), .weight_in(reg_weight_30_53), .partial_sum_in(reg_psum_30_53), .reg_activation(reg_activation_31_53), .reg_weight(reg_weight_31_53), .reg_partial_sum(reg_psum_31_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_54( .activation_in(reg_activation_31_53), .weight_in(reg_weight_30_54), .partial_sum_in(reg_psum_30_54), .reg_activation(reg_activation_31_54), .reg_weight(reg_weight_31_54), .reg_partial_sum(reg_psum_31_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_55( .activation_in(reg_activation_31_54), .weight_in(reg_weight_30_55), .partial_sum_in(reg_psum_30_55), .reg_activation(reg_activation_31_55), .reg_weight(reg_weight_31_55), .reg_partial_sum(reg_psum_31_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_56( .activation_in(reg_activation_31_55), .weight_in(reg_weight_30_56), .partial_sum_in(reg_psum_30_56), .reg_activation(reg_activation_31_56), .reg_weight(reg_weight_31_56), .reg_partial_sum(reg_psum_31_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_57( .activation_in(reg_activation_31_56), .weight_in(reg_weight_30_57), .partial_sum_in(reg_psum_30_57), .reg_activation(reg_activation_31_57), .reg_weight(reg_weight_31_57), .reg_partial_sum(reg_psum_31_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_58( .activation_in(reg_activation_31_57), .weight_in(reg_weight_30_58), .partial_sum_in(reg_psum_30_58), .reg_activation(reg_activation_31_58), .reg_weight(reg_weight_31_58), .reg_partial_sum(reg_psum_31_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_59( .activation_in(reg_activation_31_58), .weight_in(reg_weight_30_59), .partial_sum_in(reg_psum_30_59), .reg_activation(reg_activation_31_59), .reg_weight(reg_weight_31_59), .reg_partial_sum(reg_psum_31_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_60( .activation_in(reg_activation_31_59), .weight_in(reg_weight_30_60), .partial_sum_in(reg_psum_30_60), .reg_activation(reg_activation_31_60), .reg_weight(reg_weight_31_60), .reg_partial_sum(reg_psum_31_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_61( .activation_in(reg_activation_31_60), .weight_in(reg_weight_30_61), .partial_sum_in(reg_psum_30_61), .reg_activation(reg_activation_31_61), .reg_weight(reg_weight_31_61), .reg_partial_sum(reg_psum_31_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_62( .activation_in(reg_activation_31_61), .weight_in(reg_weight_30_62), .partial_sum_in(reg_psum_30_62), .reg_activation(reg_activation_31_62), .reg_weight(reg_weight_31_62), .reg_partial_sum(reg_psum_31_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_63( .activation_in(reg_activation_31_62), .weight_in(reg_weight_30_63), .partial_sum_in(reg_psum_30_63), .reg_weight(reg_weight_31_63), .reg_partial_sum(reg_psum_31_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_0( .activation_in(in_activation_32), .weight_in(reg_weight_31_0), .partial_sum_in(reg_psum_31_0), .reg_activation(reg_activation_32_0), .reg_weight(reg_weight_32_0), .reg_partial_sum(reg_psum_32_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_1( .activation_in(reg_activation_32_0), .weight_in(reg_weight_31_1), .partial_sum_in(reg_psum_31_1), .reg_activation(reg_activation_32_1), .reg_weight(reg_weight_32_1), .reg_partial_sum(reg_psum_32_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_2( .activation_in(reg_activation_32_1), .weight_in(reg_weight_31_2), .partial_sum_in(reg_psum_31_2), .reg_activation(reg_activation_32_2), .reg_weight(reg_weight_32_2), .reg_partial_sum(reg_psum_32_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_3( .activation_in(reg_activation_32_2), .weight_in(reg_weight_31_3), .partial_sum_in(reg_psum_31_3), .reg_activation(reg_activation_32_3), .reg_weight(reg_weight_32_3), .reg_partial_sum(reg_psum_32_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_4( .activation_in(reg_activation_32_3), .weight_in(reg_weight_31_4), .partial_sum_in(reg_psum_31_4), .reg_activation(reg_activation_32_4), .reg_weight(reg_weight_32_4), .reg_partial_sum(reg_psum_32_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_5( .activation_in(reg_activation_32_4), .weight_in(reg_weight_31_5), .partial_sum_in(reg_psum_31_5), .reg_activation(reg_activation_32_5), .reg_weight(reg_weight_32_5), .reg_partial_sum(reg_psum_32_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_6( .activation_in(reg_activation_32_5), .weight_in(reg_weight_31_6), .partial_sum_in(reg_psum_31_6), .reg_activation(reg_activation_32_6), .reg_weight(reg_weight_32_6), .reg_partial_sum(reg_psum_32_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_7( .activation_in(reg_activation_32_6), .weight_in(reg_weight_31_7), .partial_sum_in(reg_psum_31_7), .reg_activation(reg_activation_32_7), .reg_weight(reg_weight_32_7), .reg_partial_sum(reg_psum_32_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_8( .activation_in(reg_activation_32_7), .weight_in(reg_weight_31_8), .partial_sum_in(reg_psum_31_8), .reg_activation(reg_activation_32_8), .reg_weight(reg_weight_32_8), .reg_partial_sum(reg_psum_32_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_9( .activation_in(reg_activation_32_8), .weight_in(reg_weight_31_9), .partial_sum_in(reg_psum_31_9), .reg_activation(reg_activation_32_9), .reg_weight(reg_weight_32_9), .reg_partial_sum(reg_psum_32_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_10( .activation_in(reg_activation_32_9), .weight_in(reg_weight_31_10), .partial_sum_in(reg_psum_31_10), .reg_activation(reg_activation_32_10), .reg_weight(reg_weight_32_10), .reg_partial_sum(reg_psum_32_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_11( .activation_in(reg_activation_32_10), .weight_in(reg_weight_31_11), .partial_sum_in(reg_psum_31_11), .reg_activation(reg_activation_32_11), .reg_weight(reg_weight_32_11), .reg_partial_sum(reg_psum_32_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_12( .activation_in(reg_activation_32_11), .weight_in(reg_weight_31_12), .partial_sum_in(reg_psum_31_12), .reg_activation(reg_activation_32_12), .reg_weight(reg_weight_32_12), .reg_partial_sum(reg_psum_32_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_13( .activation_in(reg_activation_32_12), .weight_in(reg_weight_31_13), .partial_sum_in(reg_psum_31_13), .reg_activation(reg_activation_32_13), .reg_weight(reg_weight_32_13), .reg_partial_sum(reg_psum_32_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_14( .activation_in(reg_activation_32_13), .weight_in(reg_weight_31_14), .partial_sum_in(reg_psum_31_14), .reg_activation(reg_activation_32_14), .reg_weight(reg_weight_32_14), .reg_partial_sum(reg_psum_32_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_15( .activation_in(reg_activation_32_14), .weight_in(reg_weight_31_15), .partial_sum_in(reg_psum_31_15), .reg_activation(reg_activation_32_15), .reg_weight(reg_weight_32_15), .reg_partial_sum(reg_psum_32_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_16( .activation_in(reg_activation_32_15), .weight_in(reg_weight_31_16), .partial_sum_in(reg_psum_31_16), .reg_activation(reg_activation_32_16), .reg_weight(reg_weight_32_16), .reg_partial_sum(reg_psum_32_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_17( .activation_in(reg_activation_32_16), .weight_in(reg_weight_31_17), .partial_sum_in(reg_psum_31_17), .reg_activation(reg_activation_32_17), .reg_weight(reg_weight_32_17), .reg_partial_sum(reg_psum_32_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_18( .activation_in(reg_activation_32_17), .weight_in(reg_weight_31_18), .partial_sum_in(reg_psum_31_18), .reg_activation(reg_activation_32_18), .reg_weight(reg_weight_32_18), .reg_partial_sum(reg_psum_32_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_19( .activation_in(reg_activation_32_18), .weight_in(reg_weight_31_19), .partial_sum_in(reg_psum_31_19), .reg_activation(reg_activation_32_19), .reg_weight(reg_weight_32_19), .reg_partial_sum(reg_psum_32_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_20( .activation_in(reg_activation_32_19), .weight_in(reg_weight_31_20), .partial_sum_in(reg_psum_31_20), .reg_activation(reg_activation_32_20), .reg_weight(reg_weight_32_20), .reg_partial_sum(reg_psum_32_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_21( .activation_in(reg_activation_32_20), .weight_in(reg_weight_31_21), .partial_sum_in(reg_psum_31_21), .reg_activation(reg_activation_32_21), .reg_weight(reg_weight_32_21), .reg_partial_sum(reg_psum_32_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_22( .activation_in(reg_activation_32_21), .weight_in(reg_weight_31_22), .partial_sum_in(reg_psum_31_22), .reg_activation(reg_activation_32_22), .reg_weight(reg_weight_32_22), .reg_partial_sum(reg_psum_32_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_23( .activation_in(reg_activation_32_22), .weight_in(reg_weight_31_23), .partial_sum_in(reg_psum_31_23), .reg_activation(reg_activation_32_23), .reg_weight(reg_weight_32_23), .reg_partial_sum(reg_psum_32_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_24( .activation_in(reg_activation_32_23), .weight_in(reg_weight_31_24), .partial_sum_in(reg_psum_31_24), .reg_activation(reg_activation_32_24), .reg_weight(reg_weight_32_24), .reg_partial_sum(reg_psum_32_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_25( .activation_in(reg_activation_32_24), .weight_in(reg_weight_31_25), .partial_sum_in(reg_psum_31_25), .reg_activation(reg_activation_32_25), .reg_weight(reg_weight_32_25), .reg_partial_sum(reg_psum_32_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_26( .activation_in(reg_activation_32_25), .weight_in(reg_weight_31_26), .partial_sum_in(reg_psum_31_26), .reg_activation(reg_activation_32_26), .reg_weight(reg_weight_32_26), .reg_partial_sum(reg_psum_32_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_27( .activation_in(reg_activation_32_26), .weight_in(reg_weight_31_27), .partial_sum_in(reg_psum_31_27), .reg_activation(reg_activation_32_27), .reg_weight(reg_weight_32_27), .reg_partial_sum(reg_psum_32_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_28( .activation_in(reg_activation_32_27), .weight_in(reg_weight_31_28), .partial_sum_in(reg_psum_31_28), .reg_activation(reg_activation_32_28), .reg_weight(reg_weight_32_28), .reg_partial_sum(reg_psum_32_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_29( .activation_in(reg_activation_32_28), .weight_in(reg_weight_31_29), .partial_sum_in(reg_psum_31_29), .reg_activation(reg_activation_32_29), .reg_weight(reg_weight_32_29), .reg_partial_sum(reg_psum_32_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_30( .activation_in(reg_activation_32_29), .weight_in(reg_weight_31_30), .partial_sum_in(reg_psum_31_30), .reg_activation(reg_activation_32_30), .reg_weight(reg_weight_32_30), .reg_partial_sum(reg_psum_32_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_31( .activation_in(reg_activation_32_30), .weight_in(reg_weight_31_31), .partial_sum_in(reg_psum_31_31), .reg_activation(reg_activation_32_31), .reg_weight(reg_weight_32_31), .reg_partial_sum(reg_psum_32_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_32( .activation_in(reg_activation_32_31), .weight_in(reg_weight_31_32), .partial_sum_in(reg_psum_31_32), .reg_activation(reg_activation_32_32), .reg_weight(reg_weight_32_32), .reg_partial_sum(reg_psum_32_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_33( .activation_in(reg_activation_32_32), .weight_in(reg_weight_31_33), .partial_sum_in(reg_psum_31_33), .reg_activation(reg_activation_32_33), .reg_weight(reg_weight_32_33), .reg_partial_sum(reg_psum_32_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_34( .activation_in(reg_activation_32_33), .weight_in(reg_weight_31_34), .partial_sum_in(reg_psum_31_34), .reg_activation(reg_activation_32_34), .reg_weight(reg_weight_32_34), .reg_partial_sum(reg_psum_32_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_35( .activation_in(reg_activation_32_34), .weight_in(reg_weight_31_35), .partial_sum_in(reg_psum_31_35), .reg_activation(reg_activation_32_35), .reg_weight(reg_weight_32_35), .reg_partial_sum(reg_psum_32_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_36( .activation_in(reg_activation_32_35), .weight_in(reg_weight_31_36), .partial_sum_in(reg_psum_31_36), .reg_activation(reg_activation_32_36), .reg_weight(reg_weight_32_36), .reg_partial_sum(reg_psum_32_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_37( .activation_in(reg_activation_32_36), .weight_in(reg_weight_31_37), .partial_sum_in(reg_psum_31_37), .reg_activation(reg_activation_32_37), .reg_weight(reg_weight_32_37), .reg_partial_sum(reg_psum_32_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_38( .activation_in(reg_activation_32_37), .weight_in(reg_weight_31_38), .partial_sum_in(reg_psum_31_38), .reg_activation(reg_activation_32_38), .reg_weight(reg_weight_32_38), .reg_partial_sum(reg_psum_32_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_39( .activation_in(reg_activation_32_38), .weight_in(reg_weight_31_39), .partial_sum_in(reg_psum_31_39), .reg_activation(reg_activation_32_39), .reg_weight(reg_weight_32_39), .reg_partial_sum(reg_psum_32_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_40( .activation_in(reg_activation_32_39), .weight_in(reg_weight_31_40), .partial_sum_in(reg_psum_31_40), .reg_activation(reg_activation_32_40), .reg_weight(reg_weight_32_40), .reg_partial_sum(reg_psum_32_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_41( .activation_in(reg_activation_32_40), .weight_in(reg_weight_31_41), .partial_sum_in(reg_psum_31_41), .reg_activation(reg_activation_32_41), .reg_weight(reg_weight_32_41), .reg_partial_sum(reg_psum_32_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_42( .activation_in(reg_activation_32_41), .weight_in(reg_weight_31_42), .partial_sum_in(reg_psum_31_42), .reg_activation(reg_activation_32_42), .reg_weight(reg_weight_32_42), .reg_partial_sum(reg_psum_32_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_43( .activation_in(reg_activation_32_42), .weight_in(reg_weight_31_43), .partial_sum_in(reg_psum_31_43), .reg_activation(reg_activation_32_43), .reg_weight(reg_weight_32_43), .reg_partial_sum(reg_psum_32_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_44( .activation_in(reg_activation_32_43), .weight_in(reg_weight_31_44), .partial_sum_in(reg_psum_31_44), .reg_activation(reg_activation_32_44), .reg_weight(reg_weight_32_44), .reg_partial_sum(reg_psum_32_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_45( .activation_in(reg_activation_32_44), .weight_in(reg_weight_31_45), .partial_sum_in(reg_psum_31_45), .reg_activation(reg_activation_32_45), .reg_weight(reg_weight_32_45), .reg_partial_sum(reg_psum_32_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_46( .activation_in(reg_activation_32_45), .weight_in(reg_weight_31_46), .partial_sum_in(reg_psum_31_46), .reg_activation(reg_activation_32_46), .reg_weight(reg_weight_32_46), .reg_partial_sum(reg_psum_32_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_47( .activation_in(reg_activation_32_46), .weight_in(reg_weight_31_47), .partial_sum_in(reg_psum_31_47), .reg_activation(reg_activation_32_47), .reg_weight(reg_weight_32_47), .reg_partial_sum(reg_psum_32_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_48( .activation_in(reg_activation_32_47), .weight_in(reg_weight_31_48), .partial_sum_in(reg_psum_31_48), .reg_activation(reg_activation_32_48), .reg_weight(reg_weight_32_48), .reg_partial_sum(reg_psum_32_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_49( .activation_in(reg_activation_32_48), .weight_in(reg_weight_31_49), .partial_sum_in(reg_psum_31_49), .reg_activation(reg_activation_32_49), .reg_weight(reg_weight_32_49), .reg_partial_sum(reg_psum_32_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_50( .activation_in(reg_activation_32_49), .weight_in(reg_weight_31_50), .partial_sum_in(reg_psum_31_50), .reg_activation(reg_activation_32_50), .reg_weight(reg_weight_32_50), .reg_partial_sum(reg_psum_32_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_51( .activation_in(reg_activation_32_50), .weight_in(reg_weight_31_51), .partial_sum_in(reg_psum_31_51), .reg_activation(reg_activation_32_51), .reg_weight(reg_weight_32_51), .reg_partial_sum(reg_psum_32_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_52( .activation_in(reg_activation_32_51), .weight_in(reg_weight_31_52), .partial_sum_in(reg_psum_31_52), .reg_activation(reg_activation_32_52), .reg_weight(reg_weight_32_52), .reg_partial_sum(reg_psum_32_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_53( .activation_in(reg_activation_32_52), .weight_in(reg_weight_31_53), .partial_sum_in(reg_psum_31_53), .reg_activation(reg_activation_32_53), .reg_weight(reg_weight_32_53), .reg_partial_sum(reg_psum_32_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_54( .activation_in(reg_activation_32_53), .weight_in(reg_weight_31_54), .partial_sum_in(reg_psum_31_54), .reg_activation(reg_activation_32_54), .reg_weight(reg_weight_32_54), .reg_partial_sum(reg_psum_32_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_55( .activation_in(reg_activation_32_54), .weight_in(reg_weight_31_55), .partial_sum_in(reg_psum_31_55), .reg_activation(reg_activation_32_55), .reg_weight(reg_weight_32_55), .reg_partial_sum(reg_psum_32_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_56( .activation_in(reg_activation_32_55), .weight_in(reg_weight_31_56), .partial_sum_in(reg_psum_31_56), .reg_activation(reg_activation_32_56), .reg_weight(reg_weight_32_56), .reg_partial_sum(reg_psum_32_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_57( .activation_in(reg_activation_32_56), .weight_in(reg_weight_31_57), .partial_sum_in(reg_psum_31_57), .reg_activation(reg_activation_32_57), .reg_weight(reg_weight_32_57), .reg_partial_sum(reg_psum_32_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_58( .activation_in(reg_activation_32_57), .weight_in(reg_weight_31_58), .partial_sum_in(reg_psum_31_58), .reg_activation(reg_activation_32_58), .reg_weight(reg_weight_32_58), .reg_partial_sum(reg_psum_32_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_59( .activation_in(reg_activation_32_58), .weight_in(reg_weight_31_59), .partial_sum_in(reg_psum_31_59), .reg_activation(reg_activation_32_59), .reg_weight(reg_weight_32_59), .reg_partial_sum(reg_psum_32_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_60( .activation_in(reg_activation_32_59), .weight_in(reg_weight_31_60), .partial_sum_in(reg_psum_31_60), .reg_activation(reg_activation_32_60), .reg_weight(reg_weight_32_60), .reg_partial_sum(reg_psum_32_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_61( .activation_in(reg_activation_32_60), .weight_in(reg_weight_31_61), .partial_sum_in(reg_psum_31_61), .reg_activation(reg_activation_32_61), .reg_weight(reg_weight_32_61), .reg_partial_sum(reg_psum_32_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_62( .activation_in(reg_activation_32_61), .weight_in(reg_weight_31_62), .partial_sum_in(reg_psum_31_62), .reg_activation(reg_activation_32_62), .reg_weight(reg_weight_32_62), .reg_partial_sum(reg_psum_32_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U32_63( .activation_in(reg_activation_32_62), .weight_in(reg_weight_31_63), .partial_sum_in(reg_psum_31_63), .reg_weight(reg_weight_32_63), .reg_partial_sum(reg_psum_32_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_0( .activation_in(in_activation_33), .weight_in(reg_weight_32_0), .partial_sum_in(reg_psum_32_0), .reg_activation(reg_activation_33_0), .reg_weight(reg_weight_33_0), .reg_partial_sum(reg_psum_33_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_1( .activation_in(reg_activation_33_0), .weight_in(reg_weight_32_1), .partial_sum_in(reg_psum_32_1), .reg_activation(reg_activation_33_1), .reg_weight(reg_weight_33_1), .reg_partial_sum(reg_psum_33_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_2( .activation_in(reg_activation_33_1), .weight_in(reg_weight_32_2), .partial_sum_in(reg_psum_32_2), .reg_activation(reg_activation_33_2), .reg_weight(reg_weight_33_2), .reg_partial_sum(reg_psum_33_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_3( .activation_in(reg_activation_33_2), .weight_in(reg_weight_32_3), .partial_sum_in(reg_psum_32_3), .reg_activation(reg_activation_33_3), .reg_weight(reg_weight_33_3), .reg_partial_sum(reg_psum_33_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_4( .activation_in(reg_activation_33_3), .weight_in(reg_weight_32_4), .partial_sum_in(reg_psum_32_4), .reg_activation(reg_activation_33_4), .reg_weight(reg_weight_33_4), .reg_partial_sum(reg_psum_33_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_5( .activation_in(reg_activation_33_4), .weight_in(reg_weight_32_5), .partial_sum_in(reg_psum_32_5), .reg_activation(reg_activation_33_5), .reg_weight(reg_weight_33_5), .reg_partial_sum(reg_psum_33_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_6( .activation_in(reg_activation_33_5), .weight_in(reg_weight_32_6), .partial_sum_in(reg_psum_32_6), .reg_activation(reg_activation_33_6), .reg_weight(reg_weight_33_6), .reg_partial_sum(reg_psum_33_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_7( .activation_in(reg_activation_33_6), .weight_in(reg_weight_32_7), .partial_sum_in(reg_psum_32_7), .reg_activation(reg_activation_33_7), .reg_weight(reg_weight_33_7), .reg_partial_sum(reg_psum_33_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_8( .activation_in(reg_activation_33_7), .weight_in(reg_weight_32_8), .partial_sum_in(reg_psum_32_8), .reg_activation(reg_activation_33_8), .reg_weight(reg_weight_33_8), .reg_partial_sum(reg_psum_33_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_9( .activation_in(reg_activation_33_8), .weight_in(reg_weight_32_9), .partial_sum_in(reg_psum_32_9), .reg_activation(reg_activation_33_9), .reg_weight(reg_weight_33_9), .reg_partial_sum(reg_psum_33_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_10( .activation_in(reg_activation_33_9), .weight_in(reg_weight_32_10), .partial_sum_in(reg_psum_32_10), .reg_activation(reg_activation_33_10), .reg_weight(reg_weight_33_10), .reg_partial_sum(reg_psum_33_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_11( .activation_in(reg_activation_33_10), .weight_in(reg_weight_32_11), .partial_sum_in(reg_psum_32_11), .reg_activation(reg_activation_33_11), .reg_weight(reg_weight_33_11), .reg_partial_sum(reg_psum_33_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_12( .activation_in(reg_activation_33_11), .weight_in(reg_weight_32_12), .partial_sum_in(reg_psum_32_12), .reg_activation(reg_activation_33_12), .reg_weight(reg_weight_33_12), .reg_partial_sum(reg_psum_33_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_13( .activation_in(reg_activation_33_12), .weight_in(reg_weight_32_13), .partial_sum_in(reg_psum_32_13), .reg_activation(reg_activation_33_13), .reg_weight(reg_weight_33_13), .reg_partial_sum(reg_psum_33_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_14( .activation_in(reg_activation_33_13), .weight_in(reg_weight_32_14), .partial_sum_in(reg_psum_32_14), .reg_activation(reg_activation_33_14), .reg_weight(reg_weight_33_14), .reg_partial_sum(reg_psum_33_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_15( .activation_in(reg_activation_33_14), .weight_in(reg_weight_32_15), .partial_sum_in(reg_psum_32_15), .reg_activation(reg_activation_33_15), .reg_weight(reg_weight_33_15), .reg_partial_sum(reg_psum_33_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_16( .activation_in(reg_activation_33_15), .weight_in(reg_weight_32_16), .partial_sum_in(reg_psum_32_16), .reg_activation(reg_activation_33_16), .reg_weight(reg_weight_33_16), .reg_partial_sum(reg_psum_33_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_17( .activation_in(reg_activation_33_16), .weight_in(reg_weight_32_17), .partial_sum_in(reg_psum_32_17), .reg_activation(reg_activation_33_17), .reg_weight(reg_weight_33_17), .reg_partial_sum(reg_psum_33_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_18( .activation_in(reg_activation_33_17), .weight_in(reg_weight_32_18), .partial_sum_in(reg_psum_32_18), .reg_activation(reg_activation_33_18), .reg_weight(reg_weight_33_18), .reg_partial_sum(reg_psum_33_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_19( .activation_in(reg_activation_33_18), .weight_in(reg_weight_32_19), .partial_sum_in(reg_psum_32_19), .reg_activation(reg_activation_33_19), .reg_weight(reg_weight_33_19), .reg_partial_sum(reg_psum_33_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_20( .activation_in(reg_activation_33_19), .weight_in(reg_weight_32_20), .partial_sum_in(reg_psum_32_20), .reg_activation(reg_activation_33_20), .reg_weight(reg_weight_33_20), .reg_partial_sum(reg_psum_33_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_21( .activation_in(reg_activation_33_20), .weight_in(reg_weight_32_21), .partial_sum_in(reg_psum_32_21), .reg_activation(reg_activation_33_21), .reg_weight(reg_weight_33_21), .reg_partial_sum(reg_psum_33_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_22( .activation_in(reg_activation_33_21), .weight_in(reg_weight_32_22), .partial_sum_in(reg_psum_32_22), .reg_activation(reg_activation_33_22), .reg_weight(reg_weight_33_22), .reg_partial_sum(reg_psum_33_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_23( .activation_in(reg_activation_33_22), .weight_in(reg_weight_32_23), .partial_sum_in(reg_psum_32_23), .reg_activation(reg_activation_33_23), .reg_weight(reg_weight_33_23), .reg_partial_sum(reg_psum_33_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_24( .activation_in(reg_activation_33_23), .weight_in(reg_weight_32_24), .partial_sum_in(reg_psum_32_24), .reg_activation(reg_activation_33_24), .reg_weight(reg_weight_33_24), .reg_partial_sum(reg_psum_33_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_25( .activation_in(reg_activation_33_24), .weight_in(reg_weight_32_25), .partial_sum_in(reg_psum_32_25), .reg_activation(reg_activation_33_25), .reg_weight(reg_weight_33_25), .reg_partial_sum(reg_psum_33_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_26( .activation_in(reg_activation_33_25), .weight_in(reg_weight_32_26), .partial_sum_in(reg_psum_32_26), .reg_activation(reg_activation_33_26), .reg_weight(reg_weight_33_26), .reg_partial_sum(reg_psum_33_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_27( .activation_in(reg_activation_33_26), .weight_in(reg_weight_32_27), .partial_sum_in(reg_psum_32_27), .reg_activation(reg_activation_33_27), .reg_weight(reg_weight_33_27), .reg_partial_sum(reg_psum_33_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_28( .activation_in(reg_activation_33_27), .weight_in(reg_weight_32_28), .partial_sum_in(reg_psum_32_28), .reg_activation(reg_activation_33_28), .reg_weight(reg_weight_33_28), .reg_partial_sum(reg_psum_33_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_29( .activation_in(reg_activation_33_28), .weight_in(reg_weight_32_29), .partial_sum_in(reg_psum_32_29), .reg_activation(reg_activation_33_29), .reg_weight(reg_weight_33_29), .reg_partial_sum(reg_psum_33_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_30( .activation_in(reg_activation_33_29), .weight_in(reg_weight_32_30), .partial_sum_in(reg_psum_32_30), .reg_activation(reg_activation_33_30), .reg_weight(reg_weight_33_30), .reg_partial_sum(reg_psum_33_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_31( .activation_in(reg_activation_33_30), .weight_in(reg_weight_32_31), .partial_sum_in(reg_psum_32_31), .reg_activation(reg_activation_33_31), .reg_weight(reg_weight_33_31), .reg_partial_sum(reg_psum_33_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_32( .activation_in(reg_activation_33_31), .weight_in(reg_weight_32_32), .partial_sum_in(reg_psum_32_32), .reg_activation(reg_activation_33_32), .reg_weight(reg_weight_33_32), .reg_partial_sum(reg_psum_33_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_33( .activation_in(reg_activation_33_32), .weight_in(reg_weight_32_33), .partial_sum_in(reg_psum_32_33), .reg_activation(reg_activation_33_33), .reg_weight(reg_weight_33_33), .reg_partial_sum(reg_psum_33_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_34( .activation_in(reg_activation_33_33), .weight_in(reg_weight_32_34), .partial_sum_in(reg_psum_32_34), .reg_activation(reg_activation_33_34), .reg_weight(reg_weight_33_34), .reg_partial_sum(reg_psum_33_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_35( .activation_in(reg_activation_33_34), .weight_in(reg_weight_32_35), .partial_sum_in(reg_psum_32_35), .reg_activation(reg_activation_33_35), .reg_weight(reg_weight_33_35), .reg_partial_sum(reg_psum_33_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_36( .activation_in(reg_activation_33_35), .weight_in(reg_weight_32_36), .partial_sum_in(reg_psum_32_36), .reg_activation(reg_activation_33_36), .reg_weight(reg_weight_33_36), .reg_partial_sum(reg_psum_33_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_37( .activation_in(reg_activation_33_36), .weight_in(reg_weight_32_37), .partial_sum_in(reg_psum_32_37), .reg_activation(reg_activation_33_37), .reg_weight(reg_weight_33_37), .reg_partial_sum(reg_psum_33_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_38( .activation_in(reg_activation_33_37), .weight_in(reg_weight_32_38), .partial_sum_in(reg_psum_32_38), .reg_activation(reg_activation_33_38), .reg_weight(reg_weight_33_38), .reg_partial_sum(reg_psum_33_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_39( .activation_in(reg_activation_33_38), .weight_in(reg_weight_32_39), .partial_sum_in(reg_psum_32_39), .reg_activation(reg_activation_33_39), .reg_weight(reg_weight_33_39), .reg_partial_sum(reg_psum_33_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_40( .activation_in(reg_activation_33_39), .weight_in(reg_weight_32_40), .partial_sum_in(reg_psum_32_40), .reg_activation(reg_activation_33_40), .reg_weight(reg_weight_33_40), .reg_partial_sum(reg_psum_33_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_41( .activation_in(reg_activation_33_40), .weight_in(reg_weight_32_41), .partial_sum_in(reg_psum_32_41), .reg_activation(reg_activation_33_41), .reg_weight(reg_weight_33_41), .reg_partial_sum(reg_psum_33_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_42( .activation_in(reg_activation_33_41), .weight_in(reg_weight_32_42), .partial_sum_in(reg_psum_32_42), .reg_activation(reg_activation_33_42), .reg_weight(reg_weight_33_42), .reg_partial_sum(reg_psum_33_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_43( .activation_in(reg_activation_33_42), .weight_in(reg_weight_32_43), .partial_sum_in(reg_psum_32_43), .reg_activation(reg_activation_33_43), .reg_weight(reg_weight_33_43), .reg_partial_sum(reg_psum_33_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_44( .activation_in(reg_activation_33_43), .weight_in(reg_weight_32_44), .partial_sum_in(reg_psum_32_44), .reg_activation(reg_activation_33_44), .reg_weight(reg_weight_33_44), .reg_partial_sum(reg_psum_33_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_45( .activation_in(reg_activation_33_44), .weight_in(reg_weight_32_45), .partial_sum_in(reg_psum_32_45), .reg_activation(reg_activation_33_45), .reg_weight(reg_weight_33_45), .reg_partial_sum(reg_psum_33_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_46( .activation_in(reg_activation_33_45), .weight_in(reg_weight_32_46), .partial_sum_in(reg_psum_32_46), .reg_activation(reg_activation_33_46), .reg_weight(reg_weight_33_46), .reg_partial_sum(reg_psum_33_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_47( .activation_in(reg_activation_33_46), .weight_in(reg_weight_32_47), .partial_sum_in(reg_psum_32_47), .reg_activation(reg_activation_33_47), .reg_weight(reg_weight_33_47), .reg_partial_sum(reg_psum_33_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_48( .activation_in(reg_activation_33_47), .weight_in(reg_weight_32_48), .partial_sum_in(reg_psum_32_48), .reg_activation(reg_activation_33_48), .reg_weight(reg_weight_33_48), .reg_partial_sum(reg_psum_33_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_49( .activation_in(reg_activation_33_48), .weight_in(reg_weight_32_49), .partial_sum_in(reg_psum_32_49), .reg_activation(reg_activation_33_49), .reg_weight(reg_weight_33_49), .reg_partial_sum(reg_psum_33_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_50( .activation_in(reg_activation_33_49), .weight_in(reg_weight_32_50), .partial_sum_in(reg_psum_32_50), .reg_activation(reg_activation_33_50), .reg_weight(reg_weight_33_50), .reg_partial_sum(reg_psum_33_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_51( .activation_in(reg_activation_33_50), .weight_in(reg_weight_32_51), .partial_sum_in(reg_psum_32_51), .reg_activation(reg_activation_33_51), .reg_weight(reg_weight_33_51), .reg_partial_sum(reg_psum_33_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_52( .activation_in(reg_activation_33_51), .weight_in(reg_weight_32_52), .partial_sum_in(reg_psum_32_52), .reg_activation(reg_activation_33_52), .reg_weight(reg_weight_33_52), .reg_partial_sum(reg_psum_33_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_53( .activation_in(reg_activation_33_52), .weight_in(reg_weight_32_53), .partial_sum_in(reg_psum_32_53), .reg_activation(reg_activation_33_53), .reg_weight(reg_weight_33_53), .reg_partial_sum(reg_psum_33_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_54( .activation_in(reg_activation_33_53), .weight_in(reg_weight_32_54), .partial_sum_in(reg_psum_32_54), .reg_activation(reg_activation_33_54), .reg_weight(reg_weight_33_54), .reg_partial_sum(reg_psum_33_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_55( .activation_in(reg_activation_33_54), .weight_in(reg_weight_32_55), .partial_sum_in(reg_psum_32_55), .reg_activation(reg_activation_33_55), .reg_weight(reg_weight_33_55), .reg_partial_sum(reg_psum_33_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_56( .activation_in(reg_activation_33_55), .weight_in(reg_weight_32_56), .partial_sum_in(reg_psum_32_56), .reg_activation(reg_activation_33_56), .reg_weight(reg_weight_33_56), .reg_partial_sum(reg_psum_33_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_57( .activation_in(reg_activation_33_56), .weight_in(reg_weight_32_57), .partial_sum_in(reg_psum_32_57), .reg_activation(reg_activation_33_57), .reg_weight(reg_weight_33_57), .reg_partial_sum(reg_psum_33_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_58( .activation_in(reg_activation_33_57), .weight_in(reg_weight_32_58), .partial_sum_in(reg_psum_32_58), .reg_activation(reg_activation_33_58), .reg_weight(reg_weight_33_58), .reg_partial_sum(reg_psum_33_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_59( .activation_in(reg_activation_33_58), .weight_in(reg_weight_32_59), .partial_sum_in(reg_psum_32_59), .reg_activation(reg_activation_33_59), .reg_weight(reg_weight_33_59), .reg_partial_sum(reg_psum_33_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_60( .activation_in(reg_activation_33_59), .weight_in(reg_weight_32_60), .partial_sum_in(reg_psum_32_60), .reg_activation(reg_activation_33_60), .reg_weight(reg_weight_33_60), .reg_partial_sum(reg_psum_33_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_61( .activation_in(reg_activation_33_60), .weight_in(reg_weight_32_61), .partial_sum_in(reg_psum_32_61), .reg_activation(reg_activation_33_61), .reg_weight(reg_weight_33_61), .reg_partial_sum(reg_psum_33_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_62( .activation_in(reg_activation_33_61), .weight_in(reg_weight_32_62), .partial_sum_in(reg_psum_32_62), .reg_activation(reg_activation_33_62), .reg_weight(reg_weight_33_62), .reg_partial_sum(reg_psum_33_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U33_63( .activation_in(reg_activation_33_62), .weight_in(reg_weight_32_63), .partial_sum_in(reg_psum_32_63), .reg_weight(reg_weight_33_63), .reg_partial_sum(reg_psum_33_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_0( .activation_in(in_activation_34), .weight_in(reg_weight_33_0), .partial_sum_in(reg_psum_33_0), .reg_activation(reg_activation_34_0), .reg_weight(reg_weight_34_0), .reg_partial_sum(reg_psum_34_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_1( .activation_in(reg_activation_34_0), .weight_in(reg_weight_33_1), .partial_sum_in(reg_psum_33_1), .reg_activation(reg_activation_34_1), .reg_weight(reg_weight_34_1), .reg_partial_sum(reg_psum_34_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_2( .activation_in(reg_activation_34_1), .weight_in(reg_weight_33_2), .partial_sum_in(reg_psum_33_2), .reg_activation(reg_activation_34_2), .reg_weight(reg_weight_34_2), .reg_partial_sum(reg_psum_34_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_3( .activation_in(reg_activation_34_2), .weight_in(reg_weight_33_3), .partial_sum_in(reg_psum_33_3), .reg_activation(reg_activation_34_3), .reg_weight(reg_weight_34_3), .reg_partial_sum(reg_psum_34_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_4( .activation_in(reg_activation_34_3), .weight_in(reg_weight_33_4), .partial_sum_in(reg_psum_33_4), .reg_activation(reg_activation_34_4), .reg_weight(reg_weight_34_4), .reg_partial_sum(reg_psum_34_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_5( .activation_in(reg_activation_34_4), .weight_in(reg_weight_33_5), .partial_sum_in(reg_psum_33_5), .reg_activation(reg_activation_34_5), .reg_weight(reg_weight_34_5), .reg_partial_sum(reg_psum_34_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_6( .activation_in(reg_activation_34_5), .weight_in(reg_weight_33_6), .partial_sum_in(reg_psum_33_6), .reg_activation(reg_activation_34_6), .reg_weight(reg_weight_34_6), .reg_partial_sum(reg_psum_34_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_7( .activation_in(reg_activation_34_6), .weight_in(reg_weight_33_7), .partial_sum_in(reg_psum_33_7), .reg_activation(reg_activation_34_7), .reg_weight(reg_weight_34_7), .reg_partial_sum(reg_psum_34_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_8( .activation_in(reg_activation_34_7), .weight_in(reg_weight_33_8), .partial_sum_in(reg_psum_33_8), .reg_activation(reg_activation_34_8), .reg_weight(reg_weight_34_8), .reg_partial_sum(reg_psum_34_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_9( .activation_in(reg_activation_34_8), .weight_in(reg_weight_33_9), .partial_sum_in(reg_psum_33_9), .reg_activation(reg_activation_34_9), .reg_weight(reg_weight_34_9), .reg_partial_sum(reg_psum_34_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_10( .activation_in(reg_activation_34_9), .weight_in(reg_weight_33_10), .partial_sum_in(reg_psum_33_10), .reg_activation(reg_activation_34_10), .reg_weight(reg_weight_34_10), .reg_partial_sum(reg_psum_34_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_11( .activation_in(reg_activation_34_10), .weight_in(reg_weight_33_11), .partial_sum_in(reg_psum_33_11), .reg_activation(reg_activation_34_11), .reg_weight(reg_weight_34_11), .reg_partial_sum(reg_psum_34_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_12( .activation_in(reg_activation_34_11), .weight_in(reg_weight_33_12), .partial_sum_in(reg_psum_33_12), .reg_activation(reg_activation_34_12), .reg_weight(reg_weight_34_12), .reg_partial_sum(reg_psum_34_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_13( .activation_in(reg_activation_34_12), .weight_in(reg_weight_33_13), .partial_sum_in(reg_psum_33_13), .reg_activation(reg_activation_34_13), .reg_weight(reg_weight_34_13), .reg_partial_sum(reg_psum_34_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_14( .activation_in(reg_activation_34_13), .weight_in(reg_weight_33_14), .partial_sum_in(reg_psum_33_14), .reg_activation(reg_activation_34_14), .reg_weight(reg_weight_34_14), .reg_partial_sum(reg_psum_34_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_15( .activation_in(reg_activation_34_14), .weight_in(reg_weight_33_15), .partial_sum_in(reg_psum_33_15), .reg_activation(reg_activation_34_15), .reg_weight(reg_weight_34_15), .reg_partial_sum(reg_psum_34_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_16( .activation_in(reg_activation_34_15), .weight_in(reg_weight_33_16), .partial_sum_in(reg_psum_33_16), .reg_activation(reg_activation_34_16), .reg_weight(reg_weight_34_16), .reg_partial_sum(reg_psum_34_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_17( .activation_in(reg_activation_34_16), .weight_in(reg_weight_33_17), .partial_sum_in(reg_psum_33_17), .reg_activation(reg_activation_34_17), .reg_weight(reg_weight_34_17), .reg_partial_sum(reg_psum_34_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_18( .activation_in(reg_activation_34_17), .weight_in(reg_weight_33_18), .partial_sum_in(reg_psum_33_18), .reg_activation(reg_activation_34_18), .reg_weight(reg_weight_34_18), .reg_partial_sum(reg_psum_34_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_19( .activation_in(reg_activation_34_18), .weight_in(reg_weight_33_19), .partial_sum_in(reg_psum_33_19), .reg_activation(reg_activation_34_19), .reg_weight(reg_weight_34_19), .reg_partial_sum(reg_psum_34_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_20( .activation_in(reg_activation_34_19), .weight_in(reg_weight_33_20), .partial_sum_in(reg_psum_33_20), .reg_activation(reg_activation_34_20), .reg_weight(reg_weight_34_20), .reg_partial_sum(reg_psum_34_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_21( .activation_in(reg_activation_34_20), .weight_in(reg_weight_33_21), .partial_sum_in(reg_psum_33_21), .reg_activation(reg_activation_34_21), .reg_weight(reg_weight_34_21), .reg_partial_sum(reg_psum_34_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_22( .activation_in(reg_activation_34_21), .weight_in(reg_weight_33_22), .partial_sum_in(reg_psum_33_22), .reg_activation(reg_activation_34_22), .reg_weight(reg_weight_34_22), .reg_partial_sum(reg_psum_34_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_23( .activation_in(reg_activation_34_22), .weight_in(reg_weight_33_23), .partial_sum_in(reg_psum_33_23), .reg_activation(reg_activation_34_23), .reg_weight(reg_weight_34_23), .reg_partial_sum(reg_psum_34_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_24( .activation_in(reg_activation_34_23), .weight_in(reg_weight_33_24), .partial_sum_in(reg_psum_33_24), .reg_activation(reg_activation_34_24), .reg_weight(reg_weight_34_24), .reg_partial_sum(reg_psum_34_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_25( .activation_in(reg_activation_34_24), .weight_in(reg_weight_33_25), .partial_sum_in(reg_psum_33_25), .reg_activation(reg_activation_34_25), .reg_weight(reg_weight_34_25), .reg_partial_sum(reg_psum_34_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_26( .activation_in(reg_activation_34_25), .weight_in(reg_weight_33_26), .partial_sum_in(reg_psum_33_26), .reg_activation(reg_activation_34_26), .reg_weight(reg_weight_34_26), .reg_partial_sum(reg_psum_34_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_27( .activation_in(reg_activation_34_26), .weight_in(reg_weight_33_27), .partial_sum_in(reg_psum_33_27), .reg_activation(reg_activation_34_27), .reg_weight(reg_weight_34_27), .reg_partial_sum(reg_psum_34_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_28( .activation_in(reg_activation_34_27), .weight_in(reg_weight_33_28), .partial_sum_in(reg_psum_33_28), .reg_activation(reg_activation_34_28), .reg_weight(reg_weight_34_28), .reg_partial_sum(reg_psum_34_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_29( .activation_in(reg_activation_34_28), .weight_in(reg_weight_33_29), .partial_sum_in(reg_psum_33_29), .reg_activation(reg_activation_34_29), .reg_weight(reg_weight_34_29), .reg_partial_sum(reg_psum_34_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_30( .activation_in(reg_activation_34_29), .weight_in(reg_weight_33_30), .partial_sum_in(reg_psum_33_30), .reg_activation(reg_activation_34_30), .reg_weight(reg_weight_34_30), .reg_partial_sum(reg_psum_34_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_31( .activation_in(reg_activation_34_30), .weight_in(reg_weight_33_31), .partial_sum_in(reg_psum_33_31), .reg_activation(reg_activation_34_31), .reg_weight(reg_weight_34_31), .reg_partial_sum(reg_psum_34_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_32( .activation_in(reg_activation_34_31), .weight_in(reg_weight_33_32), .partial_sum_in(reg_psum_33_32), .reg_activation(reg_activation_34_32), .reg_weight(reg_weight_34_32), .reg_partial_sum(reg_psum_34_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_33( .activation_in(reg_activation_34_32), .weight_in(reg_weight_33_33), .partial_sum_in(reg_psum_33_33), .reg_activation(reg_activation_34_33), .reg_weight(reg_weight_34_33), .reg_partial_sum(reg_psum_34_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_34( .activation_in(reg_activation_34_33), .weight_in(reg_weight_33_34), .partial_sum_in(reg_psum_33_34), .reg_activation(reg_activation_34_34), .reg_weight(reg_weight_34_34), .reg_partial_sum(reg_psum_34_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_35( .activation_in(reg_activation_34_34), .weight_in(reg_weight_33_35), .partial_sum_in(reg_psum_33_35), .reg_activation(reg_activation_34_35), .reg_weight(reg_weight_34_35), .reg_partial_sum(reg_psum_34_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_36( .activation_in(reg_activation_34_35), .weight_in(reg_weight_33_36), .partial_sum_in(reg_psum_33_36), .reg_activation(reg_activation_34_36), .reg_weight(reg_weight_34_36), .reg_partial_sum(reg_psum_34_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_37( .activation_in(reg_activation_34_36), .weight_in(reg_weight_33_37), .partial_sum_in(reg_psum_33_37), .reg_activation(reg_activation_34_37), .reg_weight(reg_weight_34_37), .reg_partial_sum(reg_psum_34_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_38( .activation_in(reg_activation_34_37), .weight_in(reg_weight_33_38), .partial_sum_in(reg_psum_33_38), .reg_activation(reg_activation_34_38), .reg_weight(reg_weight_34_38), .reg_partial_sum(reg_psum_34_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_39( .activation_in(reg_activation_34_38), .weight_in(reg_weight_33_39), .partial_sum_in(reg_psum_33_39), .reg_activation(reg_activation_34_39), .reg_weight(reg_weight_34_39), .reg_partial_sum(reg_psum_34_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_40( .activation_in(reg_activation_34_39), .weight_in(reg_weight_33_40), .partial_sum_in(reg_psum_33_40), .reg_activation(reg_activation_34_40), .reg_weight(reg_weight_34_40), .reg_partial_sum(reg_psum_34_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_41( .activation_in(reg_activation_34_40), .weight_in(reg_weight_33_41), .partial_sum_in(reg_psum_33_41), .reg_activation(reg_activation_34_41), .reg_weight(reg_weight_34_41), .reg_partial_sum(reg_psum_34_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_42( .activation_in(reg_activation_34_41), .weight_in(reg_weight_33_42), .partial_sum_in(reg_psum_33_42), .reg_activation(reg_activation_34_42), .reg_weight(reg_weight_34_42), .reg_partial_sum(reg_psum_34_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_43( .activation_in(reg_activation_34_42), .weight_in(reg_weight_33_43), .partial_sum_in(reg_psum_33_43), .reg_activation(reg_activation_34_43), .reg_weight(reg_weight_34_43), .reg_partial_sum(reg_psum_34_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_44( .activation_in(reg_activation_34_43), .weight_in(reg_weight_33_44), .partial_sum_in(reg_psum_33_44), .reg_activation(reg_activation_34_44), .reg_weight(reg_weight_34_44), .reg_partial_sum(reg_psum_34_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_45( .activation_in(reg_activation_34_44), .weight_in(reg_weight_33_45), .partial_sum_in(reg_psum_33_45), .reg_activation(reg_activation_34_45), .reg_weight(reg_weight_34_45), .reg_partial_sum(reg_psum_34_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_46( .activation_in(reg_activation_34_45), .weight_in(reg_weight_33_46), .partial_sum_in(reg_psum_33_46), .reg_activation(reg_activation_34_46), .reg_weight(reg_weight_34_46), .reg_partial_sum(reg_psum_34_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_47( .activation_in(reg_activation_34_46), .weight_in(reg_weight_33_47), .partial_sum_in(reg_psum_33_47), .reg_activation(reg_activation_34_47), .reg_weight(reg_weight_34_47), .reg_partial_sum(reg_psum_34_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_48( .activation_in(reg_activation_34_47), .weight_in(reg_weight_33_48), .partial_sum_in(reg_psum_33_48), .reg_activation(reg_activation_34_48), .reg_weight(reg_weight_34_48), .reg_partial_sum(reg_psum_34_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_49( .activation_in(reg_activation_34_48), .weight_in(reg_weight_33_49), .partial_sum_in(reg_psum_33_49), .reg_activation(reg_activation_34_49), .reg_weight(reg_weight_34_49), .reg_partial_sum(reg_psum_34_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_50( .activation_in(reg_activation_34_49), .weight_in(reg_weight_33_50), .partial_sum_in(reg_psum_33_50), .reg_activation(reg_activation_34_50), .reg_weight(reg_weight_34_50), .reg_partial_sum(reg_psum_34_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_51( .activation_in(reg_activation_34_50), .weight_in(reg_weight_33_51), .partial_sum_in(reg_psum_33_51), .reg_activation(reg_activation_34_51), .reg_weight(reg_weight_34_51), .reg_partial_sum(reg_psum_34_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_52( .activation_in(reg_activation_34_51), .weight_in(reg_weight_33_52), .partial_sum_in(reg_psum_33_52), .reg_activation(reg_activation_34_52), .reg_weight(reg_weight_34_52), .reg_partial_sum(reg_psum_34_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_53( .activation_in(reg_activation_34_52), .weight_in(reg_weight_33_53), .partial_sum_in(reg_psum_33_53), .reg_activation(reg_activation_34_53), .reg_weight(reg_weight_34_53), .reg_partial_sum(reg_psum_34_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_54( .activation_in(reg_activation_34_53), .weight_in(reg_weight_33_54), .partial_sum_in(reg_psum_33_54), .reg_activation(reg_activation_34_54), .reg_weight(reg_weight_34_54), .reg_partial_sum(reg_psum_34_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_55( .activation_in(reg_activation_34_54), .weight_in(reg_weight_33_55), .partial_sum_in(reg_psum_33_55), .reg_activation(reg_activation_34_55), .reg_weight(reg_weight_34_55), .reg_partial_sum(reg_psum_34_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_56( .activation_in(reg_activation_34_55), .weight_in(reg_weight_33_56), .partial_sum_in(reg_psum_33_56), .reg_activation(reg_activation_34_56), .reg_weight(reg_weight_34_56), .reg_partial_sum(reg_psum_34_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_57( .activation_in(reg_activation_34_56), .weight_in(reg_weight_33_57), .partial_sum_in(reg_psum_33_57), .reg_activation(reg_activation_34_57), .reg_weight(reg_weight_34_57), .reg_partial_sum(reg_psum_34_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_58( .activation_in(reg_activation_34_57), .weight_in(reg_weight_33_58), .partial_sum_in(reg_psum_33_58), .reg_activation(reg_activation_34_58), .reg_weight(reg_weight_34_58), .reg_partial_sum(reg_psum_34_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_59( .activation_in(reg_activation_34_58), .weight_in(reg_weight_33_59), .partial_sum_in(reg_psum_33_59), .reg_activation(reg_activation_34_59), .reg_weight(reg_weight_34_59), .reg_partial_sum(reg_psum_34_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_60( .activation_in(reg_activation_34_59), .weight_in(reg_weight_33_60), .partial_sum_in(reg_psum_33_60), .reg_activation(reg_activation_34_60), .reg_weight(reg_weight_34_60), .reg_partial_sum(reg_psum_34_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_61( .activation_in(reg_activation_34_60), .weight_in(reg_weight_33_61), .partial_sum_in(reg_psum_33_61), .reg_activation(reg_activation_34_61), .reg_weight(reg_weight_34_61), .reg_partial_sum(reg_psum_34_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_62( .activation_in(reg_activation_34_61), .weight_in(reg_weight_33_62), .partial_sum_in(reg_psum_33_62), .reg_activation(reg_activation_34_62), .reg_weight(reg_weight_34_62), .reg_partial_sum(reg_psum_34_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U34_63( .activation_in(reg_activation_34_62), .weight_in(reg_weight_33_63), .partial_sum_in(reg_psum_33_63), .reg_weight(reg_weight_34_63), .reg_partial_sum(reg_psum_34_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_0( .activation_in(in_activation_35), .weight_in(reg_weight_34_0), .partial_sum_in(reg_psum_34_0), .reg_activation(reg_activation_35_0), .reg_weight(reg_weight_35_0), .reg_partial_sum(reg_psum_35_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_1( .activation_in(reg_activation_35_0), .weight_in(reg_weight_34_1), .partial_sum_in(reg_psum_34_1), .reg_activation(reg_activation_35_1), .reg_weight(reg_weight_35_1), .reg_partial_sum(reg_psum_35_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_2( .activation_in(reg_activation_35_1), .weight_in(reg_weight_34_2), .partial_sum_in(reg_psum_34_2), .reg_activation(reg_activation_35_2), .reg_weight(reg_weight_35_2), .reg_partial_sum(reg_psum_35_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_3( .activation_in(reg_activation_35_2), .weight_in(reg_weight_34_3), .partial_sum_in(reg_psum_34_3), .reg_activation(reg_activation_35_3), .reg_weight(reg_weight_35_3), .reg_partial_sum(reg_psum_35_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_4( .activation_in(reg_activation_35_3), .weight_in(reg_weight_34_4), .partial_sum_in(reg_psum_34_4), .reg_activation(reg_activation_35_4), .reg_weight(reg_weight_35_4), .reg_partial_sum(reg_psum_35_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_5( .activation_in(reg_activation_35_4), .weight_in(reg_weight_34_5), .partial_sum_in(reg_psum_34_5), .reg_activation(reg_activation_35_5), .reg_weight(reg_weight_35_5), .reg_partial_sum(reg_psum_35_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_6( .activation_in(reg_activation_35_5), .weight_in(reg_weight_34_6), .partial_sum_in(reg_psum_34_6), .reg_activation(reg_activation_35_6), .reg_weight(reg_weight_35_6), .reg_partial_sum(reg_psum_35_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_7( .activation_in(reg_activation_35_6), .weight_in(reg_weight_34_7), .partial_sum_in(reg_psum_34_7), .reg_activation(reg_activation_35_7), .reg_weight(reg_weight_35_7), .reg_partial_sum(reg_psum_35_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_8( .activation_in(reg_activation_35_7), .weight_in(reg_weight_34_8), .partial_sum_in(reg_psum_34_8), .reg_activation(reg_activation_35_8), .reg_weight(reg_weight_35_8), .reg_partial_sum(reg_psum_35_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_9( .activation_in(reg_activation_35_8), .weight_in(reg_weight_34_9), .partial_sum_in(reg_psum_34_9), .reg_activation(reg_activation_35_9), .reg_weight(reg_weight_35_9), .reg_partial_sum(reg_psum_35_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_10( .activation_in(reg_activation_35_9), .weight_in(reg_weight_34_10), .partial_sum_in(reg_psum_34_10), .reg_activation(reg_activation_35_10), .reg_weight(reg_weight_35_10), .reg_partial_sum(reg_psum_35_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_11( .activation_in(reg_activation_35_10), .weight_in(reg_weight_34_11), .partial_sum_in(reg_psum_34_11), .reg_activation(reg_activation_35_11), .reg_weight(reg_weight_35_11), .reg_partial_sum(reg_psum_35_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_12( .activation_in(reg_activation_35_11), .weight_in(reg_weight_34_12), .partial_sum_in(reg_psum_34_12), .reg_activation(reg_activation_35_12), .reg_weight(reg_weight_35_12), .reg_partial_sum(reg_psum_35_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_13( .activation_in(reg_activation_35_12), .weight_in(reg_weight_34_13), .partial_sum_in(reg_psum_34_13), .reg_activation(reg_activation_35_13), .reg_weight(reg_weight_35_13), .reg_partial_sum(reg_psum_35_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_14( .activation_in(reg_activation_35_13), .weight_in(reg_weight_34_14), .partial_sum_in(reg_psum_34_14), .reg_activation(reg_activation_35_14), .reg_weight(reg_weight_35_14), .reg_partial_sum(reg_psum_35_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_15( .activation_in(reg_activation_35_14), .weight_in(reg_weight_34_15), .partial_sum_in(reg_psum_34_15), .reg_activation(reg_activation_35_15), .reg_weight(reg_weight_35_15), .reg_partial_sum(reg_psum_35_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_16( .activation_in(reg_activation_35_15), .weight_in(reg_weight_34_16), .partial_sum_in(reg_psum_34_16), .reg_activation(reg_activation_35_16), .reg_weight(reg_weight_35_16), .reg_partial_sum(reg_psum_35_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_17( .activation_in(reg_activation_35_16), .weight_in(reg_weight_34_17), .partial_sum_in(reg_psum_34_17), .reg_activation(reg_activation_35_17), .reg_weight(reg_weight_35_17), .reg_partial_sum(reg_psum_35_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_18( .activation_in(reg_activation_35_17), .weight_in(reg_weight_34_18), .partial_sum_in(reg_psum_34_18), .reg_activation(reg_activation_35_18), .reg_weight(reg_weight_35_18), .reg_partial_sum(reg_psum_35_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_19( .activation_in(reg_activation_35_18), .weight_in(reg_weight_34_19), .partial_sum_in(reg_psum_34_19), .reg_activation(reg_activation_35_19), .reg_weight(reg_weight_35_19), .reg_partial_sum(reg_psum_35_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_20( .activation_in(reg_activation_35_19), .weight_in(reg_weight_34_20), .partial_sum_in(reg_psum_34_20), .reg_activation(reg_activation_35_20), .reg_weight(reg_weight_35_20), .reg_partial_sum(reg_psum_35_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_21( .activation_in(reg_activation_35_20), .weight_in(reg_weight_34_21), .partial_sum_in(reg_psum_34_21), .reg_activation(reg_activation_35_21), .reg_weight(reg_weight_35_21), .reg_partial_sum(reg_psum_35_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_22( .activation_in(reg_activation_35_21), .weight_in(reg_weight_34_22), .partial_sum_in(reg_psum_34_22), .reg_activation(reg_activation_35_22), .reg_weight(reg_weight_35_22), .reg_partial_sum(reg_psum_35_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_23( .activation_in(reg_activation_35_22), .weight_in(reg_weight_34_23), .partial_sum_in(reg_psum_34_23), .reg_activation(reg_activation_35_23), .reg_weight(reg_weight_35_23), .reg_partial_sum(reg_psum_35_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_24( .activation_in(reg_activation_35_23), .weight_in(reg_weight_34_24), .partial_sum_in(reg_psum_34_24), .reg_activation(reg_activation_35_24), .reg_weight(reg_weight_35_24), .reg_partial_sum(reg_psum_35_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_25( .activation_in(reg_activation_35_24), .weight_in(reg_weight_34_25), .partial_sum_in(reg_psum_34_25), .reg_activation(reg_activation_35_25), .reg_weight(reg_weight_35_25), .reg_partial_sum(reg_psum_35_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_26( .activation_in(reg_activation_35_25), .weight_in(reg_weight_34_26), .partial_sum_in(reg_psum_34_26), .reg_activation(reg_activation_35_26), .reg_weight(reg_weight_35_26), .reg_partial_sum(reg_psum_35_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_27( .activation_in(reg_activation_35_26), .weight_in(reg_weight_34_27), .partial_sum_in(reg_psum_34_27), .reg_activation(reg_activation_35_27), .reg_weight(reg_weight_35_27), .reg_partial_sum(reg_psum_35_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_28( .activation_in(reg_activation_35_27), .weight_in(reg_weight_34_28), .partial_sum_in(reg_psum_34_28), .reg_activation(reg_activation_35_28), .reg_weight(reg_weight_35_28), .reg_partial_sum(reg_psum_35_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_29( .activation_in(reg_activation_35_28), .weight_in(reg_weight_34_29), .partial_sum_in(reg_psum_34_29), .reg_activation(reg_activation_35_29), .reg_weight(reg_weight_35_29), .reg_partial_sum(reg_psum_35_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_30( .activation_in(reg_activation_35_29), .weight_in(reg_weight_34_30), .partial_sum_in(reg_psum_34_30), .reg_activation(reg_activation_35_30), .reg_weight(reg_weight_35_30), .reg_partial_sum(reg_psum_35_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_31( .activation_in(reg_activation_35_30), .weight_in(reg_weight_34_31), .partial_sum_in(reg_psum_34_31), .reg_activation(reg_activation_35_31), .reg_weight(reg_weight_35_31), .reg_partial_sum(reg_psum_35_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_32( .activation_in(reg_activation_35_31), .weight_in(reg_weight_34_32), .partial_sum_in(reg_psum_34_32), .reg_activation(reg_activation_35_32), .reg_weight(reg_weight_35_32), .reg_partial_sum(reg_psum_35_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_33( .activation_in(reg_activation_35_32), .weight_in(reg_weight_34_33), .partial_sum_in(reg_psum_34_33), .reg_activation(reg_activation_35_33), .reg_weight(reg_weight_35_33), .reg_partial_sum(reg_psum_35_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_34( .activation_in(reg_activation_35_33), .weight_in(reg_weight_34_34), .partial_sum_in(reg_psum_34_34), .reg_activation(reg_activation_35_34), .reg_weight(reg_weight_35_34), .reg_partial_sum(reg_psum_35_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_35( .activation_in(reg_activation_35_34), .weight_in(reg_weight_34_35), .partial_sum_in(reg_psum_34_35), .reg_activation(reg_activation_35_35), .reg_weight(reg_weight_35_35), .reg_partial_sum(reg_psum_35_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_36( .activation_in(reg_activation_35_35), .weight_in(reg_weight_34_36), .partial_sum_in(reg_psum_34_36), .reg_activation(reg_activation_35_36), .reg_weight(reg_weight_35_36), .reg_partial_sum(reg_psum_35_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_37( .activation_in(reg_activation_35_36), .weight_in(reg_weight_34_37), .partial_sum_in(reg_psum_34_37), .reg_activation(reg_activation_35_37), .reg_weight(reg_weight_35_37), .reg_partial_sum(reg_psum_35_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_38( .activation_in(reg_activation_35_37), .weight_in(reg_weight_34_38), .partial_sum_in(reg_psum_34_38), .reg_activation(reg_activation_35_38), .reg_weight(reg_weight_35_38), .reg_partial_sum(reg_psum_35_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_39( .activation_in(reg_activation_35_38), .weight_in(reg_weight_34_39), .partial_sum_in(reg_psum_34_39), .reg_activation(reg_activation_35_39), .reg_weight(reg_weight_35_39), .reg_partial_sum(reg_psum_35_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_40( .activation_in(reg_activation_35_39), .weight_in(reg_weight_34_40), .partial_sum_in(reg_psum_34_40), .reg_activation(reg_activation_35_40), .reg_weight(reg_weight_35_40), .reg_partial_sum(reg_psum_35_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_41( .activation_in(reg_activation_35_40), .weight_in(reg_weight_34_41), .partial_sum_in(reg_psum_34_41), .reg_activation(reg_activation_35_41), .reg_weight(reg_weight_35_41), .reg_partial_sum(reg_psum_35_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_42( .activation_in(reg_activation_35_41), .weight_in(reg_weight_34_42), .partial_sum_in(reg_psum_34_42), .reg_activation(reg_activation_35_42), .reg_weight(reg_weight_35_42), .reg_partial_sum(reg_psum_35_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_43( .activation_in(reg_activation_35_42), .weight_in(reg_weight_34_43), .partial_sum_in(reg_psum_34_43), .reg_activation(reg_activation_35_43), .reg_weight(reg_weight_35_43), .reg_partial_sum(reg_psum_35_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_44( .activation_in(reg_activation_35_43), .weight_in(reg_weight_34_44), .partial_sum_in(reg_psum_34_44), .reg_activation(reg_activation_35_44), .reg_weight(reg_weight_35_44), .reg_partial_sum(reg_psum_35_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_45( .activation_in(reg_activation_35_44), .weight_in(reg_weight_34_45), .partial_sum_in(reg_psum_34_45), .reg_activation(reg_activation_35_45), .reg_weight(reg_weight_35_45), .reg_partial_sum(reg_psum_35_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_46( .activation_in(reg_activation_35_45), .weight_in(reg_weight_34_46), .partial_sum_in(reg_psum_34_46), .reg_activation(reg_activation_35_46), .reg_weight(reg_weight_35_46), .reg_partial_sum(reg_psum_35_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_47( .activation_in(reg_activation_35_46), .weight_in(reg_weight_34_47), .partial_sum_in(reg_psum_34_47), .reg_activation(reg_activation_35_47), .reg_weight(reg_weight_35_47), .reg_partial_sum(reg_psum_35_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_48( .activation_in(reg_activation_35_47), .weight_in(reg_weight_34_48), .partial_sum_in(reg_psum_34_48), .reg_activation(reg_activation_35_48), .reg_weight(reg_weight_35_48), .reg_partial_sum(reg_psum_35_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_49( .activation_in(reg_activation_35_48), .weight_in(reg_weight_34_49), .partial_sum_in(reg_psum_34_49), .reg_activation(reg_activation_35_49), .reg_weight(reg_weight_35_49), .reg_partial_sum(reg_psum_35_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_50( .activation_in(reg_activation_35_49), .weight_in(reg_weight_34_50), .partial_sum_in(reg_psum_34_50), .reg_activation(reg_activation_35_50), .reg_weight(reg_weight_35_50), .reg_partial_sum(reg_psum_35_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_51( .activation_in(reg_activation_35_50), .weight_in(reg_weight_34_51), .partial_sum_in(reg_psum_34_51), .reg_activation(reg_activation_35_51), .reg_weight(reg_weight_35_51), .reg_partial_sum(reg_psum_35_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_52( .activation_in(reg_activation_35_51), .weight_in(reg_weight_34_52), .partial_sum_in(reg_psum_34_52), .reg_activation(reg_activation_35_52), .reg_weight(reg_weight_35_52), .reg_partial_sum(reg_psum_35_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_53( .activation_in(reg_activation_35_52), .weight_in(reg_weight_34_53), .partial_sum_in(reg_psum_34_53), .reg_activation(reg_activation_35_53), .reg_weight(reg_weight_35_53), .reg_partial_sum(reg_psum_35_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_54( .activation_in(reg_activation_35_53), .weight_in(reg_weight_34_54), .partial_sum_in(reg_psum_34_54), .reg_activation(reg_activation_35_54), .reg_weight(reg_weight_35_54), .reg_partial_sum(reg_psum_35_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_55( .activation_in(reg_activation_35_54), .weight_in(reg_weight_34_55), .partial_sum_in(reg_psum_34_55), .reg_activation(reg_activation_35_55), .reg_weight(reg_weight_35_55), .reg_partial_sum(reg_psum_35_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_56( .activation_in(reg_activation_35_55), .weight_in(reg_weight_34_56), .partial_sum_in(reg_psum_34_56), .reg_activation(reg_activation_35_56), .reg_weight(reg_weight_35_56), .reg_partial_sum(reg_psum_35_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_57( .activation_in(reg_activation_35_56), .weight_in(reg_weight_34_57), .partial_sum_in(reg_psum_34_57), .reg_activation(reg_activation_35_57), .reg_weight(reg_weight_35_57), .reg_partial_sum(reg_psum_35_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_58( .activation_in(reg_activation_35_57), .weight_in(reg_weight_34_58), .partial_sum_in(reg_psum_34_58), .reg_activation(reg_activation_35_58), .reg_weight(reg_weight_35_58), .reg_partial_sum(reg_psum_35_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_59( .activation_in(reg_activation_35_58), .weight_in(reg_weight_34_59), .partial_sum_in(reg_psum_34_59), .reg_activation(reg_activation_35_59), .reg_weight(reg_weight_35_59), .reg_partial_sum(reg_psum_35_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_60( .activation_in(reg_activation_35_59), .weight_in(reg_weight_34_60), .partial_sum_in(reg_psum_34_60), .reg_activation(reg_activation_35_60), .reg_weight(reg_weight_35_60), .reg_partial_sum(reg_psum_35_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_61( .activation_in(reg_activation_35_60), .weight_in(reg_weight_34_61), .partial_sum_in(reg_psum_34_61), .reg_activation(reg_activation_35_61), .reg_weight(reg_weight_35_61), .reg_partial_sum(reg_psum_35_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_62( .activation_in(reg_activation_35_61), .weight_in(reg_weight_34_62), .partial_sum_in(reg_psum_34_62), .reg_activation(reg_activation_35_62), .reg_weight(reg_weight_35_62), .reg_partial_sum(reg_psum_35_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U35_63( .activation_in(reg_activation_35_62), .weight_in(reg_weight_34_63), .partial_sum_in(reg_psum_34_63), .reg_weight(reg_weight_35_63), .reg_partial_sum(reg_psum_35_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_0( .activation_in(in_activation_36), .weight_in(reg_weight_35_0), .partial_sum_in(reg_psum_35_0), .reg_activation(reg_activation_36_0), .reg_weight(reg_weight_36_0), .reg_partial_sum(reg_psum_36_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_1( .activation_in(reg_activation_36_0), .weight_in(reg_weight_35_1), .partial_sum_in(reg_psum_35_1), .reg_activation(reg_activation_36_1), .reg_weight(reg_weight_36_1), .reg_partial_sum(reg_psum_36_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_2( .activation_in(reg_activation_36_1), .weight_in(reg_weight_35_2), .partial_sum_in(reg_psum_35_2), .reg_activation(reg_activation_36_2), .reg_weight(reg_weight_36_2), .reg_partial_sum(reg_psum_36_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_3( .activation_in(reg_activation_36_2), .weight_in(reg_weight_35_3), .partial_sum_in(reg_psum_35_3), .reg_activation(reg_activation_36_3), .reg_weight(reg_weight_36_3), .reg_partial_sum(reg_psum_36_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_4( .activation_in(reg_activation_36_3), .weight_in(reg_weight_35_4), .partial_sum_in(reg_psum_35_4), .reg_activation(reg_activation_36_4), .reg_weight(reg_weight_36_4), .reg_partial_sum(reg_psum_36_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_5( .activation_in(reg_activation_36_4), .weight_in(reg_weight_35_5), .partial_sum_in(reg_psum_35_5), .reg_activation(reg_activation_36_5), .reg_weight(reg_weight_36_5), .reg_partial_sum(reg_psum_36_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_6( .activation_in(reg_activation_36_5), .weight_in(reg_weight_35_6), .partial_sum_in(reg_psum_35_6), .reg_activation(reg_activation_36_6), .reg_weight(reg_weight_36_6), .reg_partial_sum(reg_psum_36_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_7( .activation_in(reg_activation_36_6), .weight_in(reg_weight_35_7), .partial_sum_in(reg_psum_35_7), .reg_activation(reg_activation_36_7), .reg_weight(reg_weight_36_7), .reg_partial_sum(reg_psum_36_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_8( .activation_in(reg_activation_36_7), .weight_in(reg_weight_35_8), .partial_sum_in(reg_psum_35_8), .reg_activation(reg_activation_36_8), .reg_weight(reg_weight_36_8), .reg_partial_sum(reg_psum_36_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_9( .activation_in(reg_activation_36_8), .weight_in(reg_weight_35_9), .partial_sum_in(reg_psum_35_9), .reg_activation(reg_activation_36_9), .reg_weight(reg_weight_36_9), .reg_partial_sum(reg_psum_36_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_10( .activation_in(reg_activation_36_9), .weight_in(reg_weight_35_10), .partial_sum_in(reg_psum_35_10), .reg_activation(reg_activation_36_10), .reg_weight(reg_weight_36_10), .reg_partial_sum(reg_psum_36_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_11( .activation_in(reg_activation_36_10), .weight_in(reg_weight_35_11), .partial_sum_in(reg_psum_35_11), .reg_activation(reg_activation_36_11), .reg_weight(reg_weight_36_11), .reg_partial_sum(reg_psum_36_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_12( .activation_in(reg_activation_36_11), .weight_in(reg_weight_35_12), .partial_sum_in(reg_psum_35_12), .reg_activation(reg_activation_36_12), .reg_weight(reg_weight_36_12), .reg_partial_sum(reg_psum_36_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_13( .activation_in(reg_activation_36_12), .weight_in(reg_weight_35_13), .partial_sum_in(reg_psum_35_13), .reg_activation(reg_activation_36_13), .reg_weight(reg_weight_36_13), .reg_partial_sum(reg_psum_36_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_14( .activation_in(reg_activation_36_13), .weight_in(reg_weight_35_14), .partial_sum_in(reg_psum_35_14), .reg_activation(reg_activation_36_14), .reg_weight(reg_weight_36_14), .reg_partial_sum(reg_psum_36_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_15( .activation_in(reg_activation_36_14), .weight_in(reg_weight_35_15), .partial_sum_in(reg_psum_35_15), .reg_activation(reg_activation_36_15), .reg_weight(reg_weight_36_15), .reg_partial_sum(reg_psum_36_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_16( .activation_in(reg_activation_36_15), .weight_in(reg_weight_35_16), .partial_sum_in(reg_psum_35_16), .reg_activation(reg_activation_36_16), .reg_weight(reg_weight_36_16), .reg_partial_sum(reg_psum_36_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_17( .activation_in(reg_activation_36_16), .weight_in(reg_weight_35_17), .partial_sum_in(reg_psum_35_17), .reg_activation(reg_activation_36_17), .reg_weight(reg_weight_36_17), .reg_partial_sum(reg_psum_36_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_18( .activation_in(reg_activation_36_17), .weight_in(reg_weight_35_18), .partial_sum_in(reg_psum_35_18), .reg_activation(reg_activation_36_18), .reg_weight(reg_weight_36_18), .reg_partial_sum(reg_psum_36_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_19( .activation_in(reg_activation_36_18), .weight_in(reg_weight_35_19), .partial_sum_in(reg_psum_35_19), .reg_activation(reg_activation_36_19), .reg_weight(reg_weight_36_19), .reg_partial_sum(reg_psum_36_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_20( .activation_in(reg_activation_36_19), .weight_in(reg_weight_35_20), .partial_sum_in(reg_psum_35_20), .reg_activation(reg_activation_36_20), .reg_weight(reg_weight_36_20), .reg_partial_sum(reg_psum_36_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_21( .activation_in(reg_activation_36_20), .weight_in(reg_weight_35_21), .partial_sum_in(reg_psum_35_21), .reg_activation(reg_activation_36_21), .reg_weight(reg_weight_36_21), .reg_partial_sum(reg_psum_36_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_22( .activation_in(reg_activation_36_21), .weight_in(reg_weight_35_22), .partial_sum_in(reg_psum_35_22), .reg_activation(reg_activation_36_22), .reg_weight(reg_weight_36_22), .reg_partial_sum(reg_psum_36_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_23( .activation_in(reg_activation_36_22), .weight_in(reg_weight_35_23), .partial_sum_in(reg_psum_35_23), .reg_activation(reg_activation_36_23), .reg_weight(reg_weight_36_23), .reg_partial_sum(reg_psum_36_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_24( .activation_in(reg_activation_36_23), .weight_in(reg_weight_35_24), .partial_sum_in(reg_psum_35_24), .reg_activation(reg_activation_36_24), .reg_weight(reg_weight_36_24), .reg_partial_sum(reg_psum_36_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_25( .activation_in(reg_activation_36_24), .weight_in(reg_weight_35_25), .partial_sum_in(reg_psum_35_25), .reg_activation(reg_activation_36_25), .reg_weight(reg_weight_36_25), .reg_partial_sum(reg_psum_36_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_26( .activation_in(reg_activation_36_25), .weight_in(reg_weight_35_26), .partial_sum_in(reg_psum_35_26), .reg_activation(reg_activation_36_26), .reg_weight(reg_weight_36_26), .reg_partial_sum(reg_psum_36_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_27( .activation_in(reg_activation_36_26), .weight_in(reg_weight_35_27), .partial_sum_in(reg_psum_35_27), .reg_activation(reg_activation_36_27), .reg_weight(reg_weight_36_27), .reg_partial_sum(reg_psum_36_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_28( .activation_in(reg_activation_36_27), .weight_in(reg_weight_35_28), .partial_sum_in(reg_psum_35_28), .reg_activation(reg_activation_36_28), .reg_weight(reg_weight_36_28), .reg_partial_sum(reg_psum_36_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_29( .activation_in(reg_activation_36_28), .weight_in(reg_weight_35_29), .partial_sum_in(reg_psum_35_29), .reg_activation(reg_activation_36_29), .reg_weight(reg_weight_36_29), .reg_partial_sum(reg_psum_36_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_30( .activation_in(reg_activation_36_29), .weight_in(reg_weight_35_30), .partial_sum_in(reg_psum_35_30), .reg_activation(reg_activation_36_30), .reg_weight(reg_weight_36_30), .reg_partial_sum(reg_psum_36_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_31( .activation_in(reg_activation_36_30), .weight_in(reg_weight_35_31), .partial_sum_in(reg_psum_35_31), .reg_activation(reg_activation_36_31), .reg_weight(reg_weight_36_31), .reg_partial_sum(reg_psum_36_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_32( .activation_in(reg_activation_36_31), .weight_in(reg_weight_35_32), .partial_sum_in(reg_psum_35_32), .reg_activation(reg_activation_36_32), .reg_weight(reg_weight_36_32), .reg_partial_sum(reg_psum_36_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_33( .activation_in(reg_activation_36_32), .weight_in(reg_weight_35_33), .partial_sum_in(reg_psum_35_33), .reg_activation(reg_activation_36_33), .reg_weight(reg_weight_36_33), .reg_partial_sum(reg_psum_36_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_34( .activation_in(reg_activation_36_33), .weight_in(reg_weight_35_34), .partial_sum_in(reg_psum_35_34), .reg_activation(reg_activation_36_34), .reg_weight(reg_weight_36_34), .reg_partial_sum(reg_psum_36_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_35( .activation_in(reg_activation_36_34), .weight_in(reg_weight_35_35), .partial_sum_in(reg_psum_35_35), .reg_activation(reg_activation_36_35), .reg_weight(reg_weight_36_35), .reg_partial_sum(reg_psum_36_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_36( .activation_in(reg_activation_36_35), .weight_in(reg_weight_35_36), .partial_sum_in(reg_psum_35_36), .reg_activation(reg_activation_36_36), .reg_weight(reg_weight_36_36), .reg_partial_sum(reg_psum_36_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_37( .activation_in(reg_activation_36_36), .weight_in(reg_weight_35_37), .partial_sum_in(reg_psum_35_37), .reg_activation(reg_activation_36_37), .reg_weight(reg_weight_36_37), .reg_partial_sum(reg_psum_36_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_38( .activation_in(reg_activation_36_37), .weight_in(reg_weight_35_38), .partial_sum_in(reg_psum_35_38), .reg_activation(reg_activation_36_38), .reg_weight(reg_weight_36_38), .reg_partial_sum(reg_psum_36_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_39( .activation_in(reg_activation_36_38), .weight_in(reg_weight_35_39), .partial_sum_in(reg_psum_35_39), .reg_activation(reg_activation_36_39), .reg_weight(reg_weight_36_39), .reg_partial_sum(reg_psum_36_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_40( .activation_in(reg_activation_36_39), .weight_in(reg_weight_35_40), .partial_sum_in(reg_psum_35_40), .reg_activation(reg_activation_36_40), .reg_weight(reg_weight_36_40), .reg_partial_sum(reg_psum_36_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_41( .activation_in(reg_activation_36_40), .weight_in(reg_weight_35_41), .partial_sum_in(reg_psum_35_41), .reg_activation(reg_activation_36_41), .reg_weight(reg_weight_36_41), .reg_partial_sum(reg_psum_36_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_42( .activation_in(reg_activation_36_41), .weight_in(reg_weight_35_42), .partial_sum_in(reg_psum_35_42), .reg_activation(reg_activation_36_42), .reg_weight(reg_weight_36_42), .reg_partial_sum(reg_psum_36_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_43( .activation_in(reg_activation_36_42), .weight_in(reg_weight_35_43), .partial_sum_in(reg_psum_35_43), .reg_activation(reg_activation_36_43), .reg_weight(reg_weight_36_43), .reg_partial_sum(reg_psum_36_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_44( .activation_in(reg_activation_36_43), .weight_in(reg_weight_35_44), .partial_sum_in(reg_psum_35_44), .reg_activation(reg_activation_36_44), .reg_weight(reg_weight_36_44), .reg_partial_sum(reg_psum_36_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_45( .activation_in(reg_activation_36_44), .weight_in(reg_weight_35_45), .partial_sum_in(reg_psum_35_45), .reg_activation(reg_activation_36_45), .reg_weight(reg_weight_36_45), .reg_partial_sum(reg_psum_36_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_46( .activation_in(reg_activation_36_45), .weight_in(reg_weight_35_46), .partial_sum_in(reg_psum_35_46), .reg_activation(reg_activation_36_46), .reg_weight(reg_weight_36_46), .reg_partial_sum(reg_psum_36_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_47( .activation_in(reg_activation_36_46), .weight_in(reg_weight_35_47), .partial_sum_in(reg_psum_35_47), .reg_activation(reg_activation_36_47), .reg_weight(reg_weight_36_47), .reg_partial_sum(reg_psum_36_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_48( .activation_in(reg_activation_36_47), .weight_in(reg_weight_35_48), .partial_sum_in(reg_psum_35_48), .reg_activation(reg_activation_36_48), .reg_weight(reg_weight_36_48), .reg_partial_sum(reg_psum_36_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_49( .activation_in(reg_activation_36_48), .weight_in(reg_weight_35_49), .partial_sum_in(reg_psum_35_49), .reg_activation(reg_activation_36_49), .reg_weight(reg_weight_36_49), .reg_partial_sum(reg_psum_36_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_50( .activation_in(reg_activation_36_49), .weight_in(reg_weight_35_50), .partial_sum_in(reg_psum_35_50), .reg_activation(reg_activation_36_50), .reg_weight(reg_weight_36_50), .reg_partial_sum(reg_psum_36_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_51( .activation_in(reg_activation_36_50), .weight_in(reg_weight_35_51), .partial_sum_in(reg_psum_35_51), .reg_activation(reg_activation_36_51), .reg_weight(reg_weight_36_51), .reg_partial_sum(reg_psum_36_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_52( .activation_in(reg_activation_36_51), .weight_in(reg_weight_35_52), .partial_sum_in(reg_psum_35_52), .reg_activation(reg_activation_36_52), .reg_weight(reg_weight_36_52), .reg_partial_sum(reg_psum_36_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_53( .activation_in(reg_activation_36_52), .weight_in(reg_weight_35_53), .partial_sum_in(reg_psum_35_53), .reg_activation(reg_activation_36_53), .reg_weight(reg_weight_36_53), .reg_partial_sum(reg_psum_36_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_54( .activation_in(reg_activation_36_53), .weight_in(reg_weight_35_54), .partial_sum_in(reg_psum_35_54), .reg_activation(reg_activation_36_54), .reg_weight(reg_weight_36_54), .reg_partial_sum(reg_psum_36_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_55( .activation_in(reg_activation_36_54), .weight_in(reg_weight_35_55), .partial_sum_in(reg_psum_35_55), .reg_activation(reg_activation_36_55), .reg_weight(reg_weight_36_55), .reg_partial_sum(reg_psum_36_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_56( .activation_in(reg_activation_36_55), .weight_in(reg_weight_35_56), .partial_sum_in(reg_psum_35_56), .reg_activation(reg_activation_36_56), .reg_weight(reg_weight_36_56), .reg_partial_sum(reg_psum_36_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_57( .activation_in(reg_activation_36_56), .weight_in(reg_weight_35_57), .partial_sum_in(reg_psum_35_57), .reg_activation(reg_activation_36_57), .reg_weight(reg_weight_36_57), .reg_partial_sum(reg_psum_36_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_58( .activation_in(reg_activation_36_57), .weight_in(reg_weight_35_58), .partial_sum_in(reg_psum_35_58), .reg_activation(reg_activation_36_58), .reg_weight(reg_weight_36_58), .reg_partial_sum(reg_psum_36_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_59( .activation_in(reg_activation_36_58), .weight_in(reg_weight_35_59), .partial_sum_in(reg_psum_35_59), .reg_activation(reg_activation_36_59), .reg_weight(reg_weight_36_59), .reg_partial_sum(reg_psum_36_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_60( .activation_in(reg_activation_36_59), .weight_in(reg_weight_35_60), .partial_sum_in(reg_psum_35_60), .reg_activation(reg_activation_36_60), .reg_weight(reg_weight_36_60), .reg_partial_sum(reg_psum_36_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_61( .activation_in(reg_activation_36_60), .weight_in(reg_weight_35_61), .partial_sum_in(reg_psum_35_61), .reg_activation(reg_activation_36_61), .reg_weight(reg_weight_36_61), .reg_partial_sum(reg_psum_36_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_62( .activation_in(reg_activation_36_61), .weight_in(reg_weight_35_62), .partial_sum_in(reg_psum_35_62), .reg_activation(reg_activation_36_62), .reg_weight(reg_weight_36_62), .reg_partial_sum(reg_psum_36_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U36_63( .activation_in(reg_activation_36_62), .weight_in(reg_weight_35_63), .partial_sum_in(reg_psum_35_63), .reg_weight(reg_weight_36_63), .reg_partial_sum(reg_psum_36_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_0( .activation_in(in_activation_37), .weight_in(reg_weight_36_0), .partial_sum_in(reg_psum_36_0), .reg_activation(reg_activation_37_0), .reg_weight(reg_weight_37_0), .reg_partial_sum(reg_psum_37_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_1( .activation_in(reg_activation_37_0), .weight_in(reg_weight_36_1), .partial_sum_in(reg_psum_36_1), .reg_activation(reg_activation_37_1), .reg_weight(reg_weight_37_1), .reg_partial_sum(reg_psum_37_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_2( .activation_in(reg_activation_37_1), .weight_in(reg_weight_36_2), .partial_sum_in(reg_psum_36_2), .reg_activation(reg_activation_37_2), .reg_weight(reg_weight_37_2), .reg_partial_sum(reg_psum_37_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_3( .activation_in(reg_activation_37_2), .weight_in(reg_weight_36_3), .partial_sum_in(reg_psum_36_3), .reg_activation(reg_activation_37_3), .reg_weight(reg_weight_37_3), .reg_partial_sum(reg_psum_37_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_4( .activation_in(reg_activation_37_3), .weight_in(reg_weight_36_4), .partial_sum_in(reg_psum_36_4), .reg_activation(reg_activation_37_4), .reg_weight(reg_weight_37_4), .reg_partial_sum(reg_psum_37_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_5( .activation_in(reg_activation_37_4), .weight_in(reg_weight_36_5), .partial_sum_in(reg_psum_36_5), .reg_activation(reg_activation_37_5), .reg_weight(reg_weight_37_5), .reg_partial_sum(reg_psum_37_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_6( .activation_in(reg_activation_37_5), .weight_in(reg_weight_36_6), .partial_sum_in(reg_psum_36_6), .reg_activation(reg_activation_37_6), .reg_weight(reg_weight_37_6), .reg_partial_sum(reg_psum_37_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_7( .activation_in(reg_activation_37_6), .weight_in(reg_weight_36_7), .partial_sum_in(reg_psum_36_7), .reg_activation(reg_activation_37_7), .reg_weight(reg_weight_37_7), .reg_partial_sum(reg_psum_37_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_8( .activation_in(reg_activation_37_7), .weight_in(reg_weight_36_8), .partial_sum_in(reg_psum_36_8), .reg_activation(reg_activation_37_8), .reg_weight(reg_weight_37_8), .reg_partial_sum(reg_psum_37_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_9( .activation_in(reg_activation_37_8), .weight_in(reg_weight_36_9), .partial_sum_in(reg_psum_36_9), .reg_activation(reg_activation_37_9), .reg_weight(reg_weight_37_9), .reg_partial_sum(reg_psum_37_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_10( .activation_in(reg_activation_37_9), .weight_in(reg_weight_36_10), .partial_sum_in(reg_psum_36_10), .reg_activation(reg_activation_37_10), .reg_weight(reg_weight_37_10), .reg_partial_sum(reg_psum_37_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_11( .activation_in(reg_activation_37_10), .weight_in(reg_weight_36_11), .partial_sum_in(reg_psum_36_11), .reg_activation(reg_activation_37_11), .reg_weight(reg_weight_37_11), .reg_partial_sum(reg_psum_37_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_12( .activation_in(reg_activation_37_11), .weight_in(reg_weight_36_12), .partial_sum_in(reg_psum_36_12), .reg_activation(reg_activation_37_12), .reg_weight(reg_weight_37_12), .reg_partial_sum(reg_psum_37_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_13( .activation_in(reg_activation_37_12), .weight_in(reg_weight_36_13), .partial_sum_in(reg_psum_36_13), .reg_activation(reg_activation_37_13), .reg_weight(reg_weight_37_13), .reg_partial_sum(reg_psum_37_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_14( .activation_in(reg_activation_37_13), .weight_in(reg_weight_36_14), .partial_sum_in(reg_psum_36_14), .reg_activation(reg_activation_37_14), .reg_weight(reg_weight_37_14), .reg_partial_sum(reg_psum_37_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_15( .activation_in(reg_activation_37_14), .weight_in(reg_weight_36_15), .partial_sum_in(reg_psum_36_15), .reg_activation(reg_activation_37_15), .reg_weight(reg_weight_37_15), .reg_partial_sum(reg_psum_37_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_16( .activation_in(reg_activation_37_15), .weight_in(reg_weight_36_16), .partial_sum_in(reg_psum_36_16), .reg_activation(reg_activation_37_16), .reg_weight(reg_weight_37_16), .reg_partial_sum(reg_psum_37_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_17( .activation_in(reg_activation_37_16), .weight_in(reg_weight_36_17), .partial_sum_in(reg_psum_36_17), .reg_activation(reg_activation_37_17), .reg_weight(reg_weight_37_17), .reg_partial_sum(reg_psum_37_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_18( .activation_in(reg_activation_37_17), .weight_in(reg_weight_36_18), .partial_sum_in(reg_psum_36_18), .reg_activation(reg_activation_37_18), .reg_weight(reg_weight_37_18), .reg_partial_sum(reg_psum_37_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_19( .activation_in(reg_activation_37_18), .weight_in(reg_weight_36_19), .partial_sum_in(reg_psum_36_19), .reg_activation(reg_activation_37_19), .reg_weight(reg_weight_37_19), .reg_partial_sum(reg_psum_37_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_20( .activation_in(reg_activation_37_19), .weight_in(reg_weight_36_20), .partial_sum_in(reg_psum_36_20), .reg_activation(reg_activation_37_20), .reg_weight(reg_weight_37_20), .reg_partial_sum(reg_psum_37_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_21( .activation_in(reg_activation_37_20), .weight_in(reg_weight_36_21), .partial_sum_in(reg_psum_36_21), .reg_activation(reg_activation_37_21), .reg_weight(reg_weight_37_21), .reg_partial_sum(reg_psum_37_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_22( .activation_in(reg_activation_37_21), .weight_in(reg_weight_36_22), .partial_sum_in(reg_psum_36_22), .reg_activation(reg_activation_37_22), .reg_weight(reg_weight_37_22), .reg_partial_sum(reg_psum_37_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_23( .activation_in(reg_activation_37_22), .weight_in(reg_weight_36_23), .partial_sum_in(reg_psum_36_23), .reg_activation(reg_activation_37_23), .reg_weight(reg_weight_37_23), .reg_partial_sum(reg_psum_37_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_24( .activation_in(reg_activation_37_23), .weight_in(reg_weight_36_24), .partial_sum_in(reg_psum_36_24), .reg_activation(reg_activation_37_24), .reg_weight(reg_weight_37_24), .reg_partial_sum(reg_psum_37_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_25( .activation_in(reg_activation_37_24), .weight_in(reg_weight_36_25), .partial_sum_in(reg_psum_36_25), .reg_activation(reg_activation_37_25), .reg_weight(reg_weight_37_25), .reg_partial_sum(reg_psum_37_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_26( .activation_in(reg_activation_37_25), .weight_in(reg_weight_36_26), .partial_sum_in(reg_psum_36_26), .reg_activation(reg_activation_37_26), .reg_weight(reg_weight_37_26), .reg_partial_sum(reg_psum_37_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_27( .activation_in(reg_activation_37_26), .weight_in(reg_weight_36_27), .partial_sum_in(reg_psum_36_27), .reg_activation(reg_activation_37_27), .reg_weight(reg_weight_37_27), .reg_partial_sum(reg_psum_37_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_28( .activation_in(reg_activation_37_27), .weight_in(reg_weight_36_28), .partial_sum_in(reg_psum_36_28), .reg_activation(reg_activation_37_28), .reg_weight(reg_weight_37_28), .reg_partial_sum(reg_psum_37_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_29( .activation_in(reg_activation_37_28), .weight_in(reg_weight_36_29), .partial_sum_in(reg_psum_36_29), .reg_activation(reg_activation_37_29), .reg_weight(reg_weight_37_29), .reg_partial_sum(reg_psum_37_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_30( .activation_in(reg_activation_37_29), .weight_in(reg_weight_36_30), .partial_sum_in(reg_psum_36_30), .reg_activation(reg_activation_37_30), .reg_weight(reg_weight_37_30), .reg_partial_sum(reg_psum_37_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_31( .activation_in(reg_activation_37_30), .weight_in(reg_weight_36_31), .partial_sum_in(reg_psum_36_31), .reg_activation(reg_activation_37_31), .reg_weight(reg_weight_37_31), .reg_partial_sum(reg_psum_37_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_32( .activation_in(reg_activation_37_31), .weight_in(reg_weight_36_32), .partial_sum_in(reg_psum_36_32), .reg_activation(reg_activation_37_32), .reg_weight(reg_weight_37_32), .reg_partial_sum(reg_psum_37_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_33( .activation_in(reg_activation_37_32), .weight_in(reg_weight_36_33), .partial_sum_in(reg_psum_36_33), .reg_activation(reg_activation_37_33), .reg_weight(reg_weight_37_33), .reg_partial_sum(reg_psum_37_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_34( .activation_in(reg_activation_37_33), .weight_in(reg_weight_36_34), .partial_sum_in(reg_psum_36_34), .reg_activation(reg_activation_37_34), .reg_weight(reg_weight_37_34), .reg_partial_sum(reg_psum_37_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_35( .activation_in(reg_activation_37_34), .weight_in(reg_weight_36_35), .partial_sum_in(reg_psum_36_35), .reg_activation(reg_activation_37_35), .reg_weight(reg_weight_37_35), .reg_partial_sum(reg_psum_37_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_36( .activation_in(reg_activation_37_35), .weight_in(reg_weight_36_36), .partial_sum_in(reg_psum_36_36), .reg_activation(reg_activation_37_36), .reg_weight(reg_weight_37_36), .reg_partial_sum(reg_psum_37_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_37( .activation_in(reg_activation_37_36), .weight_in(reg_weight_36_37), .partial_sum_in(reg_psum_36_37), .reg_activation(reg_activation_37_37), .reg_weight(reg_weight_37_37), .reg_partial_sum(reg_psum_37_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_38( .activation_in(reg_activation_37_37), .weight_in(reg_weight_36_38), .partial_sum_in(reg_psum_36_38), .reg_activation(reg_activation_37_38), .reg_weight(reg_weight_37_38), .reg_partial_sum(reg_psum_37_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_39( .activation_in(reg_activation_37_38), .weight_in(reg_weight_36_39), .partial_sum_in(reg_psum_36_39), .reg_activation(reg_activation_37_39), .reg_weight(reg_weight_37_39), .reg_partial_sum(reg_psum_37_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_40( .activation_in(reg_activation_37_39), .weight_in(reg_weight_36_40), .partial_sum_in(reg_psum_36_40), .reg_activation(reg_activation_37_40), .reg_weight(reg_weight_37_40), .reg_partial_sum(reg_psum_37_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_41( .activation_in(reg_activation_37_40), .weight_in(reg_weight_36_41), .partial_sum_in(reg_psum_36_41), .reg_activation(reg_activation_37_41), .reg_weight(reg_weight_37_41), .reg_partial_sum(reg_psum_37_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_42( .activation_in(reg_activation_37_41), .weight_in(reg_weight_36_42), .partial_sum_in(reg_psum_36_42), .reg_activation(reg_activation_37_42), .reg_weight(reg_weight_37_42), .reg_partial_sum(reg_psum_37_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_43( .activation_in(reg_activation_37_42), .weight_in(reg_weight_36_43), .partial_sum_in(reg_psum_36_43), .reg_activation(reg_activation_37_43), .reg_weight(reg_weight_37_43), .reg_partial_sum(reg_psum_37_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_44( .activation_in(reg_activation_37_43), .weight_in(reg_weight_36_44), .partial_sum_in(reg_psum_36_44), .reg_activation(reg_activation_37_44), .reg_weight(reg_weight_37_44), .reg_partial_sum(reg_psum_37_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_45( .activation_in(reg_activation_37_44), .weight_in(reg_weight_36_45), .partial_sum_in(reg_psum_36_45), .reg_activation(reg_activation_37_45), .reg_weight(reg_weight_37_45), .reg_partial_sum(reg_psum_37_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_46( .activation_in(reg_activation_37_45), .weight_in(reg_weight_36_46), .partial_sum_in(reg_psum_36_46), .reg_activation(reg_activation_37_46), .reg_weight(reg_weight_37_46), .reg_partial_sum(reg_psum_37_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_47( .activation_in(reg_activation_37_46), .weight_in(reg_weight_36_47), .partial_sum_in(reg_psum_36_47), .reg_activation(reg_activation_37_47), .reg_weight(reg_weight_37_47), .reg_partial_sum(reg_psum_37_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_48( .activation_in(reg_activation_37_47), .weight_in(reg_weight_36_48), .partial_sum_in(reg_psum_36_48), .reg_activation(reg_activation_37_48), .reg_weight(reg_weight_37_48), .reg_partial_sum(reg_psum_37_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_49( .activation_in(reg_activation_37_48), .weight_in(reg_weight_36_49), .partial_sum_in(reg_psum_36_49), .reg_activation(reg_activation_37_49), .reg_weight(reg_weight_37_49), .reg_partial_sum(reg_psum_37_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_50( .activation_in(reg_activation_37_49), .weight_in(reg_weight_36_50), .partial_sum_in(reg_psum_36_50), .reg_activation(reg_activation_37_50), .reg_weight(reg_weight_37_50), .reg_partial_sum(reg_psum_37_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_51( .activation_in(reg_activation_37_50), .weight_in(reg_weight_36_51), .partial_sum_in(reg_psum_36_51), .reg_activation(reg_activation_37_51), .reg_weight(reg_weight_37_51), .reg_partial_sum(reg_psum_37_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_52( .activation_in(reg_activation_37_51), .weight_in(reg_weight_36_52), .partial_sum_in(reg_psum_36_52), .reg_activation(reg_activation_37_52), .reg_weight(reg_weight_37_52), .reg_partial_sum(reg_psum_37_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_53( .activation_in(reg_activation_37_52), .weight_in(reg_weight_36_53), .partial_sum_in(reg_psum_36_53), .reg_activation(reg_activation_37_53), .reg_weight(reg_weight_37_53), .reg_partial_sum(reg_psum_37_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_54( .activation_in(reg_activation_37_53), .weight_in(reg_weight_36_54), .partial_sum_in(reg_psum_36_54), .reg_activation(reg_activation_37_54), .reg_weight(reg_weight_37_54), .reg_partial_sum(reg_psum_37_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_55( .activation_in(reg_activation_37_54), .weight_in(reg_weight_36_55), .partial_sum_in(reg_psum_36_55), .reg_activation(reg_activation_37_55), .reg_weight(reg_weight_37_55), .reg_partial_sum(reg_psum_37_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_56( .activation_in(reg_activation_37_55), .weight_in(reg_weight_36_56), .partial_sum_in(reg_psum_36_56), .reg_activation(reg_activation_37_56), .reg_weight(reg_weight_37_56), .reg_partial_sum(reg_psum_37_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_57( .activation_in(reg_activation_37_56), .weight_in(reg_weight_36_57), .partial_sum_in(reg_psum_36_57), .reg_activation(reg_activation_37_57), .reg_weight(reg_weight_37_57), .reg_partial_sum(reg_psum_37_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_58( .activation_in(reg_activation_37_57), .weight_in(reg_weight_36_58), .partial_sum_in(reg_psum_36_58), .reg_activation(reg_activation_37_58), .reg_weight(reg_weight_37_58), .reg_partial_sum(reg_psum_37_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_59( .activation_in(reg_activation_37_58), .weight_in(reg_weight_36_59), .partial_sum_in(reg_psum_36_59), .reg_activation(reg_activation_37_59), .reg_weight(reg_weight_37_59), .reg_partial_sum(reg_psum_37_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_60( .activation_in(reg_activation_37_59), .weight_in(reg_weight_36_60), .partial_sum_in(reg_psum_36_60), .reg_activation(reg_activation_37_60), .reg_weight(reg_weight_37_60), .reg_partial_sum(reg_psum_37_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_61( .activation_in(reg_activation_37_60), .weight_in(reg_weight_36_61), .partial_sum_in(reg_psum_36_61), .reg_activation(reg_activation_37_61), .reg_weight(reg_weight_37_61), .reg_partial_sum(reg_psum_37_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_62( .activation_in(reg_activation_37_61), .weight_in(reg_weight_36_62), .partial_sum_in(reg_psum_36_62), .reg_activation(reg_activation_37_62), .reg_weight(reg_weight_37_62), .reg_partial_sum(reg_psum_37_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U37_63( .activation_in(reg_activation_37_62), .weight_in(reg_weight_36_63), .partial_sum_in(reg_psum_36_63), .reg_weight(reg_weight_37_63), .reg_partial_sum(reg_psum_37_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_0( .activation_in(in_activation_38), .weight_in(reg_weight_37_0), .partial_sum_in(reg_psum_37_0), .reg_activation(reg_activation_38_0), .reg_weight(reg_weight_38_0), .reg_partial_sum(reg_psum_38_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_1( .activation_in(reg_activation_38_0), .weight_in(reg_weight_37_1), .partial_sum_in(reg_psum_37_1), .reg_activation(reg_activation_38_1), .reg_weight(reg_weight_38_1), .reg_partial_sum(reg_psum_38_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_2( .activation_in(reg_activation_38_1), .weight_in(reg_weight_37_2), .partial_sum_in(reg_psum_37_2), .reg_activation(reg_activation_38_2), .reg_weight(reg_weight_38_2), .reg_partial_sum(reg_psum_38_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_3( .activation_in(reg_activation_38_2), .weight_in(reg_weight_37_3), .partial_sum_in(reg_psum_37_3), .reg_activation(reg_activation_38_3), .reg_weight(reg_weight_38_3), .reg_partial_sum(reg_psum_38_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_4( .activation_in(reg_activation_38_3), .weight_in(reg_weight_37_4), .partial_sum_in(reg_psum_37_4), .reg_activation(reg_activation_38_4), .reg_weight(reg_weight_38_4), .reg_partial_sum(reg_psum_38_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_5( .activation_in(reg_activation_38_4), .weight_in(reg_weight_37_5), .partial_sum_in(reg_psum_37_5), .reg_activation(reg_activation_38_5), .reg_weight(reg_weight_38_5), .reg_partial_sum(reg_psum_38_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_6( .activation_in(reg_activation_38_5), .weight_in(reg_weight_37_6), .partial_sum_in(reg_psum_37_6), .reg_activation(reg_activation_38_6), .reg_weight(reg_weight_38_6), .reg_partial_sum(reg_psum_38_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_7( .activation_in(reg_activation_38_6), .weight_in(reg_weight_37_7), .partial_sum_in(reg_psum_37_7), .reg_activation(reg_activation_38_7), .reg_weight(reg_weight_38_7), .reg_partial_sum(reg_psum_38_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_8( .activation_in(reg_activation_38_7), .weight_in(reg_weight_37_8), .partial_sum_in(reg_psum_37_8), .reg_activation(reg_activation_38_8), .reg_weight(reg_weight_38_8), .reg_partial_sum(reg_psum_38_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_9( .activation_in(reg_activation_38_8), .weight_in(reg_weight_37_9), .partial_sum_in(reg_psum_37_9), .reg_activation(reg_activation_38_9), .reg_weight(reg_weight_38_9), .reg_partial_sum(reg_psum_38_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_10( .activation_in(reg_activation_38_9), .weight_in(reg_weight_37_10), .partial_sum_in(reg_psum_37_10), .reg_activation(reg_activation_38_10), .reg_weight(reg_weight_38_10), .reg_partial_sum(reg_psum_38_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_11( .activation_in(reg_activation_38_10), .weight_in(reg_weight_37_11), .partial_sum_in(reg_psum_37_11), .reg_activation(reg_activation_38_11), .reg_weight(reg_weight_38_11), .reg_partial_sum(reg_psum_38_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_12( .activation_in(reg_activation_38_11), .weight_in(reg_weight_37_12), .partial_sum_in(reg_psum_37_12), .reg_activation(reg_activation_38_12), .reg_weight(reg_weight_38_12), .reg_partial_sum(reg_psum_38_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_13( .activation_in(reg_activation_38_12), .weight_in(reg_weight_37_13), .partial_sum_in(reg_psum_37_13), .reg_activation(reg_activation_38_13), .reg_weight(reg_weight_38_13), .reg_partial_sum(reg_psum_38_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_14( .activation_in(reg_activation_38_13), .weight_in(reg_weight_37_14), .partial_sum_in(reg_psum_37_14), .reg_activation(reg_activation_38_14), .reg_weight(reg_weight_38_14), .reg_partial_sum(reg_psum_38_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_15( .activation_in(reg_activation_38_14), .weight_in(reg_weight_37_15), .partial_sum_in(reg_psum_37_15), .reg_activation(reg_activation_38_15), .reg_weight(reg_weight_38_15), .reg_partial_sum(reg_psum_38_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_16( .activation_in(reg_activation_38_15), .weight_in(reg_weight_37_16), .partial_sum_in(reg_psum_37_16), .reg_activation(reg_activation_38_16), .reg_weight(reg_weight_38_16), .reg_partial_sum(reg_psum_38_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_17( .activation_in(reg_activation_38_16), .weight_in(reg_weight_37_17), .partial_sum_in(reg_psum_37_17), .reg_activation(reg_activation_38_17), .reg_weight(reg_weight_38_17), .reg_partial_sum(reg_psum_38_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_18( .activation_in(reg_activation_38_17), .weight_in(reg_weight_37_18), .partial_sum_in(reg_psum_37_18), .reg_activation(reg_activation_38_18), .reg_weight(reg_weight_38_18), .reg_partial_sum(reg_psum_38_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_19( .activation_in(reg_activation_38_18), .weight_in(reg_weight_37_19), .partial_sum_in(reg_psum_37_19), .reg_activation(reg_activation_38_19), .reg_weight(reg_weight_38_19), .reg_partial_sum(reg_psum_38_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_20( .activation_in(reg_activation_38_19), .weight_in(reg_weight_37_20), .partial_sum_in(reg_psum_37_20), .reg_activation(reg_activation_38_20), .reg_weight(reg_weight_38_20), .reg_partial_sum(reg_psum_38_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_21( .activation_in(reg_activation_38_20), .weight_in(reg_weight_37_21), .partial_sum_in(reg_psum_37_21), .reg_activation(reg_activation_38_21), .reg_weight(reg_weight_38_21), .reg_partial_sum(reg_psum_38_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_22( .activation_in(reg_activation_38_21), .weight_in(reg_weight_37_22), .partial_sum_in(reg_psum_37_22), .reg_activation(reg_activation_38_22), .reg_weight(reg_weight_38_22), .reg_partial_sum(reg_psum_38_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_23( .activation_in(reg_activation_38_22), .weight_in(reg_weight_37_23), .partial_sum_in(reg_psum_37_23), .reg_activation(reg_activation_38_23), .reg_weight(reg_weight_38_23), .reg_partial_sum(reg_psum_38_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_24( .activation_in(reg_activation_38_23), .weight_in(reg_weight_37_24), .partial_sum_in(reg_psum_37_24), .reg_activation(reg_activation_38_24), .reg_weight(reg_weight_38_24), .reg_partial_sum(reg_psum_38_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_25( .activation_in(reg_activation_38_24), .weight_in(reg_weight_37_25), .partial_sum_in(reg_psum_37_25), .reg_activation(reg_activation_38_25), .reg_weight(reg_weight_38_25), .reg_partial_sum(reg_psum_38_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_26( .activation_in(reg_activation_38_25), .weight_in(reg_weight_37_26), .partial_sum_in(reg_psum_37_26), .reg_activation(reg_activation_38_26), .reg_weight(reg_weight_38_26), .reg_partial_sum(reg_psum_38_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_27( .activation_in(reg_activation_38_26), .weight_in(reg_weight_37_27), .partial_sum_in(reg_psum_37_27), .reg_activation(reg_activation_38_27), .reg_weight(reg_weight_38_27), .reg_partial_sum(reg_psum_38_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_28( .activation_in(reg_activation_38_27), .weight_in(reg_weight_37_28), .partial_sum_in(reg_psum_37_28), .reg_activation(reg_activation_38_28), .reg_weight(reg_weight_38_28), .reg_partial_sum(reg_psum_38_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_29( .activation_in(reg_activation_38_28), .weight_in(reg_weight_37_29), .partial_sum_in(reg_psum_37_29), .reg_activation(reg_activation_38_29), .reg_weight(reg_weight_38_29), .reg_partial_sum(reg_psum_38_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_30( .activation_in(reg_activation_38_29), .weight_in(reg_weight_37_30), .partial_sum_in(reg_psum_37_30), .reg_activation(reg_activation_38_30), .reg_weight(reg_weight_38_30), .reg_partial_sum(reg_psum_38_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_31( .activation_in(reg_activation_38_30), .weight_in(reg_weight_37_31), .partial_sum_in(reg_psum_37_31), .reg_activation(reg_activation_38_31), .reg_weight(reg_weight_38_31), .reg_partial_sum(reg_psum_38_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_32( .activation_in(reg_activation_38_31), .weight_in(reg_weight_37_32), .partial_sum_in(reg_psum_37_32), .reg_activation(reg_activation_38_32), .reg_weight(reg_weight_38_32), .reg_partial_sum(reg_psum_38_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_33( .activation_in(reg_activation_38_32), .weight_in(reg_weight_37_33), .partial_sum_in(reg_psum_37_33), .reg_activation(reg_activation_38_33), .reg_weight(reg_weight_38_33), .reg_partial_sum(reg_psum_38_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_34( .activation_in(reg_activation_38_33), .weight_in(reg_weight_37_34), .partial_sum_in(reg_psum_37_34), .reg_activation(reg_activation_38_34), .reg_weight(reg_weight_38_34), .reg_partial_sum(reg_psum_38_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_35( .activation_in(reg_activation_38_34), .weight_in(reg_weight_37_35), .partial_sum_in(reg_psum_37_35), .reg_activation(reg_activation_38_35), .reg_weight(reg_weight_38_35), .reg_partial_sum(reg_psum_38_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_36( .activation_in(reg_activation_38_35), .weight_in(reg_weight_37_36), .partial_sum_in(reg_psum_37_36), .reg_activation(reg_activation_38_36), .reg_weight(reg_weight_38_36), .reg_partial_sum(reg_psum_38_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_37( .activation_in(reg_activation_38_36), .weight_in(reg_weight_37_37), .partial_sum_in(reg_psum_37_37), .reg_activation(reg_activation_38_37), .reg_weight(reg_weight_38_37), .reg_partial_sum(reg_psum_38_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_38( .activation_in(reg_activation_38_37), .weight_in(reg_weight_37_38), .partial_sum_in(reg_psum_37_38), .reg_activation(reg_activation_38_38), .reg_weight(reg_weight_38_38), .reg_partial_sum(reg_psum_38_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_39( .activation_in(reg_activation_38_38), .weight_in(reg_weight_37_39), .partial_sum_in(reg_psum_37_39), .reg_activation(reg_activation_38_39), .reg_weight(reg_weight_38_39), .reg_partial_sum(reg_psum_38_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_40( .activation_in(reg_activation_38_39), .weight_in(reg_weight_37_40), .partial_sum_in(reg_psum_37_40), .reg_activation(reg_activation_38_40), .reg_weight(reg_weight_38_40), .reg_partial_sum(reg_psum_38_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_41( .activation_in(reg_activation_38_40), .weight_in(reg_weight_37_41), .partial_sum_in(reg_psum_37_41), .reg_activation(reg_activation_38_41), .reg_weight(reg_weight_38_41), .reg_partial_sum(reg_psum_38_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_42( .activation_in(reg_activation_38_41), .weight_in(reg_weight_37_42), .partial_sum_in(reg_psum_37_42), .reg_activation(reg_activation_38_42), .reg_weight(reg_weight_38_42), .reg_partial_sum(reg_psum_38_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_43( .activation_in(reg_activation_38_42), .weight_in(reg_weight_37_43), .partial_sum_in(reg_psum_37_43), .reg_activation(reg_activation_38_43), .reg_weight(reg_weight_38_43), .reg_partial_sum(reg_psum_38_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_44( .activation_in(reg_activation_38_43), .weight_in(reg_weight_37_44), .partial_sum_in(reg_psum_37_44), .reg_activation(reg_activation_38_44), .reg_weight(reg_weight_38_44), .reg_partial_sum(reg_psum_38_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_45( .activation_in(reg_activation_38_44), .weight_in(reg_weight_37_45), .partial_sum_in(reg_psum_37_45), .reg_activation(reg_activation_38_45), .reg_weight(reg_weight_38_45), .reg_partial_sum(reg_psum_38_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_46( .activation_in(reg_activation_38_45), .weight_in(reg_weight_37_46), .partial_sum_in(reg_psum_37_46), .reg_activation(reg_activation_38_46), .reg_weight(reg_weight_38_46), .reg_partial_sum(reg_psum_38_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_47( .activation_in(reg_activation_38_46), .weight_in(reg_weight_37_47), .partial_sum_in(reg_psum_37_47), .reg_activation(reg_activation_38_47), .reg_weight(reg_weight_38_47), .reg_partial_sum(reg_psum_38_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_48( .activation_in(reg_activation_38_47), .weight_in(reg_weight_37_48), .partial_sum_in(reg_psum_37_48), .reg_activation(reg_activation_38_48), .reg_weight(reg_weight_38_48), .reg_partial_sum(reg_psum_38_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_49( .activation_in(reg_activation_38_48), .weight_in(reg_weight_37_49), .partial_sum_in(reg_psum_37_49), .reg_activation(reg_activation_38_49), .reg_weight(reg_weight_38_49), .reg_partial_sum(reg_psum_38_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_50( .activation_in(reg_activation_38_49), .weight_in(reg_weight_37_50), .partial_sum_in(reg_psum_37_50), .reg_activation(reg_activation_38_50), .reg_weight(reg_weight_38_50), .reg_partial_sum(reg_psum_38_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_51( .activation_in(reg_activation_38_50), .weight_in(reg_weight_37_51), .partial_sum_in(reg_psum_37_51), .reg_activation(reg_activation_38_51), .reg_weight(reg_weight_38_51), .reg_partial_sum(reg_psum_38_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_52( .activation_in(reg_activation_38_51), .weight_in(reg_weight_37_52), .partial_sum_in(reg_psum_37_52), .reg_activation(reg_activation_38_52), .reg_weight(reg_weight_38_52), .reg_partial_sum(reg_psum_38_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_53( .activation_in(reg_activation_38_52), .weight_in(reg_weight_37_53), .partial_sum_in(reg_psum_37_53), .reg_activation(reg_activation_38_53), .reg_weight(reg_weight_38_53), .reg_partial_sum(reg_psum_38_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_54( .activation_in(reg_activation_38_53), .weight_in(reg_weight_37_54), .partial_sum_in(reg_psum_37_54), .reg_activation(reg_activation_38_54), .reg_weight(reg_weight_38_54), .reg_partial_sum(reg_psum_38_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_55( .activation_in(reg_activation_38_54), .weight_in(reg_weight_37_55), .partial_sum_in(reg_psum_37_55), .reg_activation(reg_activation_38_55), .reg_weight(reg_weight_38_55), .reg_partial_sum(reg_psum_38_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_56( .activation_in(reg_activation_38_55), .weight_in(reg_weight_37_56), .partial_sum_in(reg_psum_37_56), .reg_activation(reg_activation_38_56), .reg_weight(reg_weight_38_56), .reg_partial_sum(reg_psum_38_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_57( .activation_in(reg_activation_38_56), .weight_in(reg_weight_37_57), .partial_sum_in(reg_psum_37_57), .reg_activation(reg_activation_38_57), .reg_weight(reg_weight_38_57), .reg_partial_sum(reg_psum_38_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_58( .activation_in(reg_activation_38_57), .weight_in(reg_weight_37_58), .partial_sum_in(reg_psum_37_58), .reg_activation(reg_activation_38_58), .reg_weight(reg_weight_38_58), .reg_partial_sum(reg_psum_38_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_59( .activation_in(reg_activation_38_58), .weight_in(reg_weight_37_59), .partial_sum_in(reg_psum_37_59), .reg_activation(reg_activation_38_59), .reg_weight(reg_weight_38_59), .reg_partial_sum(reg_psum_38_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_60( .activation_in(reg_activation_38_59), .weight_in(reg_weight_37_60), .partial_sum_in(reg_psum_37_60), .reg_activation(reg_activation_38_60), .reg_weight(reg_weight_38_60), .reg_partial_sum(reg_psum_38_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_61( .activation_in(reg_activation_38_60), .weight_in(reg_weight_37_61), .partial_sum_in(reg_psum_37_61), .reg_activation(reg_activation_38_61), .reg_weight(reg_weight_38_61), .reg_partial_sum(reg_psum_38_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_62( .activation_in(reg_activation_38_61), .weight_in(reg_weight_37_62), .partial_sum_in(reg_psum_37_62), .reg_activation(reg_activation_38_62), .reg_weight(reg_weight_38_62), .reg_partial_sum(reg_psum_38_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U38_63( .activation_in(reg_activation_38_62), .weight_in(reg_weight_37_63), .partial_sum_in(reg_psum_37_63), .reg_weight(reg_weight_38_63), .reg_partial_sum(reg_psum_38_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_0( .activation_in(in_activation_39), .weight_in(reg_weight_38_0), .partial_sum_in(reg_psum_38_0), .reg_activation(reg_activation_39_0), .reg_weight(reg_weight_39_0), .reg_partial_sum(reg_psum_39_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_1( .activation_in(reg_activation_39_0), .weight_in(reg_weight_38_1), .partial_sum_in(reg_psum_38_1), .reg_activation(reg_activation_39_1), .reg_weight(reg_weight_39_1), .reg_partial_sum(reg_psum_39_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_2( .activation_in(reg_activation_39_1), .weight_in(reg_weight_38_2), .partial_sum_in(reg_psum_38_2), .reg_activation(reg_activation_39_2), .reg_weight(reg_weight_39_2), .reg_partial_sum(reg_psum_39_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_3( .activation_in(reg_activation_39_2), .weight_in(reg_weight_38_3), .partial_sum_in(reg_psum_38_3), .reg_activation(reg_activation_39_3), .reg_weight(reg_weight_39_3), .reg_partial_sum(reg_psum_39_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_4( .activation_in(reg_activation_39_3), .weight_in(reg_weight_38_4), .partial_sum_in(reg_psum_38_4), .reg_activation(reg_activation_39_4), .reg_weight(reg_weight_39_4), .reg_partial_sum(reg_psum_39_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_5( .activation_in(reg_activation_39_4), .weight_in(reg_weight_38_5), .partial_sum_in(reg_psum_38_5), .reg_activation(reg_activation_39_5), .reg_weight(reg_weight_39_5), .reg_partial_sum(reg_psum_39_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_6( .activation_in(reg_activation_39_5), .weight_in(reg_weight_38_6), .partial_sum_in(reg_psum_38_6), .reg_activation(reg_activation_39_6), .reg_weight(reg_weight_39_6), .reg_partial_sum(reg_psum_39_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_7( .activation_in(reg_activation_39_6), .weight_in(reg_weight_38_7), .partial_sum_in(reg_psum_38_7), .reg_activation(reg_activation_39_7), .reg_weight(reg_weight_39_7), .reg_partial_sum(reg_psum_39_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_8( .activation_in(reg_activation_39_7), .weight_in(reg_weight_38_8), .partial_sum_in(reg_psum_38_8), .reg_activation(reg_activation_39_8), .reg_weight(reg_weight_39_8), .reg_partial_sum(reg_psum_39_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_9( .activation_in(reg_activation_39_8), .weight_in(reg_weight_38_9), .partial_sum_in(reg_psum_38_9), .reg_activation(reg_activation_39_9), .reg_weight(reg_weight_39_9), .reg_partial_sum(reg_psum_39_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_10( .activation_in(reg_activation_39_9), .weight_in(reg_weight_38_10), .partial_sum_in(reg_psum_38_10), .reg_activation(reg_activation_39_10), .reg_weight(reg_weight_39_10), .reg_partial_sum(reg_psum_39_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_11( .activation_in(reg_activation_39_10), .weight_in(reg_weight_38_11), .partial_sum_in(reg_psum_38_11), .reg_activation(reg_activation_39_11), .reg_weight(reg_weight_39_11), .reg_partial_sum(reg_psum_39_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_12( .activation_in(reg_activation_39_11), .weight_in(reg_weight_38_12), .partial_sum_in(reg_psum_38_12), .reg_activation(reg_activation_39_12), .reg_weight(reg_weight_39_12), .reg_partial_sum(reg_psum_39_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_13( .activation_in(reg_activation_39_12), .weight_in(reg_weight_38_13), .partial_sum_in(reg_psum_38_13), .reg_activation(reg_activation_39_13), .reg_weight(reg_weight_39_13), .reg_partial_sum(reg_psum_39_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_14( .activation_in(reg_activation_39_13), .weight_in(reg_weight_38_14), .partial_sum_in(reg_psum_38_14), .reg_activation(reg_activation_39_14), .reg_weight(reg_weight_39_14), .reg_partial_sum(reg_psum_39_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_15( .activation_in(reg_activation_39_14), .weight_in(reg_weight_38_15), .partial_sum_in(reg_psum_38_15), .reg_activation(reg_activation_39_15), .reg_weight(reg_weight_39_15), .reg_partial_sum(reg_psum_39_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_16( .activation_in(reg_activation_39_15), .weight_in(reg_weight_38_16), .partial_sum_in(reg_psum_38_16), .reg_activation(reg_activation_39_16), .reg_weight(reg_weight_39_16), .reg_partial_sum(reg_psum_39_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_17( .activation_in(reg_activation_39_16), .weight_in(reg_weight_38_17), .partial_sum_in(reg_psum_38_17), .reg_activation(reg_activation_39_17), .reg_weight(reg_weight_39_17), .reg_partial_sum(reg_psum_39_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_18( .activation_in(reg_activation_39_17), .weight_in(reg_weight_38_18), .partial_sum_in(reg_psum_38_18), .reg_activation(reg_activation_39_18), .reg_weight(reg_weight_39_18), .reg_partial_sum(reg_psum_39_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_19( .activation_in(reg_activation_39_18), .weight_in(reg_weight_38_19), .partial_sum_in(reg_psum_38_19), .reg_activation(reg_activation_39_19), .reg_weight(reg_weight_39_19), .reg_partial_sum(reg_psum_39_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_20( .activation_in(reg_activation_39_19), .weight_in(reg_weight_38_20), .partial_sum_in(reg_psum_38_20), .reg_activation(reg_activation_39_20), .reg_weight(reg_weight_39_20), .reg_partial_sum(reg_psum_39_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_21( .activation_in(reg_activation_39_20), .weight_in(reg_weight_38_21), .partial_sum_in(reg_psum_38_21), .reg_activation(reg_activation_39_21), .reg_weight(reg_weight_39_21), .reg_partial_sum(reg_psum_39_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_22( .activation_in(reg_activation_39_21), .weight_in(reg_weight_38_22), .partial_sum_in(reg_psum_38_22), .reg_activation(reg_activation_39_22), .reg_weight(reg_weight_39_22), .reg_partial_sum(reg_psum_39_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_23( .activation_in(reg_activation_39_22), .weight_in(reg_weight_38_23), .partial_sum_in(reg_psum_38_23), .reg_activation(reg_activation_39_23), .reg_weight(reg_weight_39_23), .reg_partial_sum(reg_psum_39_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_24( .activation_in(reg_activation_39_23), .weight_in(reg_weight_38_24), .partial_sum_in(reg_psum_38_24), .reg_activation(reg_activation_39_24), .reg_weight(reg_weight_39_24), .reg_partial_sum(reg_psum_39_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_25( .activation_in(reg_activation_39_24), .weight_in(reg_weight_38_25), .partial_sum_in(reg_psum_38_25), .reg_activation(reg_activation_39_25), .reg_weight(reg_weight_39_25), .reg_partial_sum(reg_psum_39_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_26( .activation_in(reg_activation_39_25), .weight_in(reg_weight_38_26), .partial_sum_in(reg_psum_38_26), .reg_activation(reg_activation_39_26), .reg_weight(reg_weight_39_26), .reg_partial_sum(reg_psum_39_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_27( .activation_in(reg_activation_39_26), .weight_in(reg_weight_38_27), .partial_sum_in(reg_psum_38_27), .reg_activation(reg_activation_39_27), .reg_weight(reg_weight_39_27), .reg_partial_sum(reg_psum_39_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_28( .activation_in(reg_activation_39_27), .weight_in(reg_weight_38_28), .partial_sum_in(reg_psum_38_28), .reg_activation(reg_activation_39_28), .reg_weight(reg_weight_39_28), .reg_partial_sum(reg_psum_39_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_29( .activation_in(reg_activation_39_28), .weight_in(reg_weight_38_29), .partial_sum_in(reg_psum_38_29), .reg_activation(reg_activation_39_29), .reg_weight(reg_weight_39_29), .reg_partial_sum(reg_psum_39_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_30( .activation_in(reg_activation_39_29), .weight_in(reg_weight_38_30), .partial_sum_in(reg_psum_38_30), .reg_activation(reg_activation_39_30), .reg_weight(reg_weight_39_30), .reg_partial_sum(reg_psum_39_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_31( .activation_in(reg_activation_39_30), .weight_in(reg_weight_38_31), .partial_sum_in(reg_psum_38_31), .reg_activation(reg_activation_39_31), .reg_weight(reg_weight_39_31), .reg_partial_sum(reg_psum_39_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_32( .activation_in(reg_activation_39_31), .weight_in(reg_weight_38_32), .partial_sum_in(reg_psum_38_32), .reg_activation(reg_activation_39_32), .reg_weight(reg_weight_39_32), .reg_partial_sum(reg_psum_39_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_33( .activation_in(reg_activation_39_32), .weight_in(reg_weight_38_33), .partial_sum_in(reg_psum_38_33), .reg_activation(reg_activation_39_33), .reg_weight(reg_weight_39_33), .reg_partial_sum(reg_psum_39_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_34( .activation_in(reg_activation_39_33), .weight_in(reg_weight_38_34), .partial_sum_in(reg_psum_38_34), .reg_activation(reg_activation_39_34), .reg_weight(reg_weight_39_34), .reg_partial_sum(reg_psum_39_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_35( .activation_in(reg_activation_39_34), .weight_in(reg_weight_38_35), .partial_sum_in(reg_psum_38_35), .reg_activation(reg_activation_39_35), .reg_weight(reg_weight_39_35), .reg_partial_sum(reg_psum_39_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_36( .activation_in(reg_activation_39_35), .weight_in(reg_weight_38_36), .partial_sum_in(reg_psum_38_36), .reg_activation(reg_activation_39_36), .reg_weight(reg_weight_39_36), .reg_partial_sum(reg_psum_39_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_37( .activation_in(reg_activation_39_36), .weight_in(reg_weight_38_37), .partial_sum_in(reg_psum_38_37), .reg_activation(reg_activation_39_37), .reg_weight(reg_weight_39_37), .reg_partial_sum(reg_psum_39_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_38( .activation_in(reg_activation_39_37), .weight_in(reg_weight_38_38), .partial_sum_in(reg_psum_38_38), .reg_activation(reg_activation_39_38), .reg_weight(reg_weight_39_38), .reg_partial_sum(reg_psum_39_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_39( .activation_in(reg_activation_39_38), .weight_in(reg_weight_38_39), .partial_sum_in(reg_psum_38_39), .reg_activation(reg_activation_39_39), .reg_weight(reg_weight_39_39), .reg_partial_sum(reg_psum_39_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_40( .activation_in(reg_activation_39_39), .weight_in(reg_weight_38_40), .partial_sum_in(reg_psum_38_40), .reg_activation(reg_activation_39_40), .reg_weight(reg_weight_39_40), .reg_partial_sum(reg_psum_39_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_41( .activation_in(reg_activation_39_40), .weight_in(reg_weight_38_41), .partial_sum_in(reg_psum_38_41), .reg_activation(reg_activation_39_41), .reg_weight(reg_weight_39_41), .reg_partial_sum(reg_psum_39_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_42( .activation_in(reg_activation_39_41), .weight_in(reg_weight_38_42), .partial_sum_in(reg_psum_38_42), .reg_activation(reg_activation_39_42), .reg_weight(reg_weight_39_42), .reg_partial_sum(reg_psum_39_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_43( .activation_in(reg_activation_39_42), .weight_in(reg_weight_38_43), .partial_sum_in(reg_psum_38_43), .reg_activation(reg_activation_39_43), .reg_weight(reg_weight_39_43), .reg_partial_sum(reg_psum_39_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_44( .activation_in(reg_activation_39_43), .weight_in(reg_weight_38_44), .partial_sum_in(reg_psum_38_44), .reg_activation(reg_activation_39_44), .reg_weight(reg_weight_39_44), .reg_partial_sum(reg_psum_39_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_45( .activation_in(reg_activation_39_44), .weight_in(reg_weight_38_45), .partial_sum_in(reg_psum_38_45), .reg_activation(reg_activation_39_45), .reg_weight(reg_weight_39_45), .reg_partial_sum(reg_psum_39_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_46( .activation_in(reg_activation_39_45), .weight_in(reg_weight_38_46), .partial_sum_in(reg_psum_38_46), .reg_activation(reg_activation_39_46), .reg_weight(reg_weight_39_46), .reg_partial_sum(reg_psum_39_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_47( .activation_in(reg_activation_39_46), .weight_in(reg_weight_38_47), .partial_sum_in(reg_psum_38_47), .reg_activation(reg_activation_39_47), .reg_weight(reg_weight_39_47), .reg_partial_sum(reg_psum_39_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_48( .activation_in(reg_activation_39_47), .weight_in(reg_weight_38_48), .partial_sum_in(reg_psum_38_48), .reg_activation(reg_activation_39_48), .reg_weight(reg_weight_39_48), .reg_partial_sum(reg_psum_39_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_49( .activation_in(reg_activation_39_48), .weight_in(reg_weight_38_49), .partial_sum_in(reg_psum_38_49), .reg_activation(reg_activation_39_49), .reg_weight(reg_weight_39_49), .reg_partial_sum(reg_psum_39_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_50( .activation_in(reg_activation_39_49), .weight_in(reg_weight_38_50), .partial_sum_in(reg_psum_38_50), .reg_activation(reg_activation_39_50), .reg_weight(reg_weight_39_50), .reg_partial_sum(reg_psum_39_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_51( .activation_in(reg_activation_39_50), .weight_in(reg_weight_38_51), .partial_sum_in(reg_psum_38_51), .reg_activation(reg_activation_39_51), .reg_weight(reg_weight_39_51), .reg_partial_sum(reg_psum_39_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_52( .activation_in(reg_activation_39_51), .weight_in(reg_weight_38_52), .partial_sum_in(reg_psum_38_52), .reg_activation(reg_activation_39_52), .reg_weight(reg_weight_39_52), .reg_partial_sum(reg_psum_39_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_53( .activation_in(reg_activation_39_52), .weight_in(reg_weight_38_53), .partial_sum_in(reg_psum_38_53), .reg_activation(reg_activation_39_53), .reg_weight(reg_weight_39_53), .reg_partial_sum(reg_psum_39_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_54( .activation_in(reg_activation_39_53), .weight_in(reg_weight_38_54), .partial_sum_in(reg_psum_38_54), .reg_activation(reg_activation_39_54), .reg_weight(reg_weight_39_54), .reg_partial_sum(reg_psum_39_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_55( .activation_in(reg_activation_39_54), .weight_in(reg_weight_38_55), .partial_sum_in(reg_psum_38_55), .reg_activation(reg_activation_39_55), .reg_weight(reg_weight_39_55), .reg_partial_sum(reg_psum_39_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_56( .activation_in(reg_activation_39_55), .weight_in(reg_weight_38_56), .partial_sum_in(reg_psum_38_56), .reg_activation(reg_activation_39_56), .reg_weight(reg_weight_39_56), .reg_partial_sum(reg_psum_39_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_57( .activation_in(reg_activation_39_56), .weight_in(reg_weight_38_57), .partial_sum_in(reg_psum_38_57), .reg_activation(reg_activation_39_57), .reg_weight(reg_weight_39_57), .reg_partial_sum(reg_psum_39_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_58( .activation_in(reg_activation_39_57), .weight_in(reg_weight_38_58), .partial_sum_in(reg_psum_38_58), .reg_activation(reg_activation_39_58), .reg_weight(reg_weight_39_58), .reg_partial_sum(reg_psum_39_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_59( .activation_in(reg_activation_39_58), .weight_in(reg_weight_38_59), .partial_sum_in(reg_psum_38_59), .reg_activation(reg_activation_39_59), .reg_weight(reg_weight_39_59), .reg_partial_sum(reg_psum_39_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_60( .activation_in(reg_activation_39_59), .weight_in(reg_weight_38_60), .partial_sum_in(reg_psum_38_60), .reg_activation(reg_activation_39_60), .reg_weight(reg_weight_39_60), .reg_partial_sum(reg_psum_39_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_61( .activation_in(reg_activation_39_60), .weight_in(reg_weight_38_61), .partial_sum_in(reg_psum_38_61), .reg_activation(reg_activation_39_61), .reg_weight(reg_weight_39_61), .reg_partial_sum(reg_psum_39_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_62( .activation_in(reg_activation_39_61), .weight_in(reg_weight_38_62), .partial_sum_in(reg_psum_38_62), .reg_activation(reg_activation_39_62), .reg_weight(reg_weight_39_62), .reg_partial_sum(reg_psum_39_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U39_63( .activation_in(reg_activation_39_62), .weight_in(reg_weight_38_63), .partial_sum_in(reg_psum_38_63), .reg_weight(reg_weight_39_63), .reg_partial_sum(reg_psum_39_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_0( .activation_in(in_activation_40), .weight_in(reg_weight_39_0), .partial_sum_in(reg_psum_39_0), .reg_activation(reg_activation_40_0), .reg_weight(reg_weight_40_0), .reg_partial_sum(reg_psum_40_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_1( .activation_in(reg_activation_40_0), .weight_in(reg_weight_39_1), .partial_sum_in(reg_psum_39_1), .reg_activation(reg_activation_40_1), .reg_weight(reg_weight_40_1), .reg_partial_sum(reg_psum_40_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_2( .activation_in(reg_activation_40_1), .weight_in(reg_weight_39_2), .partial_sum_in(reg_psum_39_2), .reg_activation(reg_activation_40_2), .reg_weight(reg_weight_40_2), .reg_partial_sum(reg_psum_40_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_3( .activation_in(reg_activation_40_2), .weight_in(reg_weight_39_3), .partial_sum_in(reg_psum_39_3), .reg_activation(reg_activation_40_3), .reg_weight(reg_weight_40_3), .reg_partial_sum(reg_psum_40_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_4( .activation_in(reg_activation_40_3), .weight_in(reg_weight_39_4), .partial_sum_in(reg_psum_39_4), .reg_activation(reg_activation_40_4), .reg_weight(reg_weight_40_4), .reg_partial_sum(reg_psum_40_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_5( .activation_in(reg_activation_40_4), .weight_in(reg_weight_39_5), .partial_sum_in(reg_psum_39_5), .reg_activation(reg_activation_40_5), .reg_weight(reg_weight_40_5), .reg_partial_sum(reg_psum_40_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_6( .activation_in(reg_activation_40_5), .weight_in(reg_weight_39_6), .partial_sum_in(reg_psum_39_6), .reg_activation(reg_activation_40_6), .reg_weight(reg_weight_40_6), .reg_partial_sum(reg_psum_40_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_7( .activation_in(reg_activation_40_6), .weight_in(reg_weight_39_7), .partial_sum_in(reg_psum_39_7), .reg_activation(reg_activation_40_7), .reg_weight(reg_weight_40_7), .reg_partial_sum(reg_psum_40_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_8( .activation_in(reg_activation_40_7), .weight_in(reg_weight_39_8), .partial_sum_in(reg_psum_39_8), .reg_activation(reg_activation_40_8), .reg_weight(reg_weight_40_8), .reg_partial_sum(reg_psum_40_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_9( .activation_in(reg_activation_40_8), .weight_in(reg_weight_39_9), .partial_sum_in(reg_psum_39_9), .reg_activation(reg_activation_40_9), .reg_weight(reg_weight_40_9), .reg_partial_sum(reg_psum_40_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_10( .activation_in(reg_activation_40_9), .weight_in(reg_weight_39_10), .partial_sum_in(reg_psum_39_10), .reg_activation(reg_activation_40_10), .reg_weight(reg_weight_40_10), .reg_partial_sum(reg_psum_40_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_11( .activation_in(reg_activation_40_10), .weight_in(reg_weight_39_11), .partial_sum_in(reg_psum_39_11), .reg_activation(reg_activation_40_11), .reg_weight(reg_weight_40_11), .reg_partial_sum(reg_psum_40_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_12( .activation_in(reg_activation_40_11), .weight_in(reg_weight_39_12), .partial_sum_in(reg_psum_39_12), .reg_activation(reg_activation_40_12), .reg_weight(reg_weight_40_12), .reg_partial_sum(reg_psum_40_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_13( .activation_in(reg_activation_40_12), .weight_in(reg_weight_39_13), .partial_sum_in(reg_psum_39_13), .reg_activation(reg_activation_40_13), .reg_weight(reg_weight_40_13), .reg_partial_sum(reg_psum_40_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_14( .activation_in(reg_activation_40_13), .weight_in(reg_weight_39_14), .partial_sum_in(reg_psum_39_14), .reg_activation(reg_activation_40_14), .reg_weight(reg_weight_40_14), .reg_partial_sum(reg_psum_40_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_15( .activation_in(reg_activation_40_14), .weight_in(reg_weight_39_15), .partial_sum_in(reg_psum_39_15), .reg_activation(reg_activation_40_15), .reg_weight(reg_weight_40_15), .reg_partial_sum(reg_psum_40_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_16( .activation_in(reg_activation_40_15), .weight_in(reg_weight_39_16), .partial_sum_in(reg_psum_39_16), .reg_activation(reg_activation_40_16), .reg_weight(reg_weight_40_16), .reg_partial_sum(reg_psum_40_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_17( .activation_in(reg_activation_40_16), .weight_in(reg_weight_39_17), .partial_sum_in(reg_psum_39_17), .reg_activation(reg_activation_40_17), .reg_weight(reg_weight_40_17), .reg_partial_sum(reg_psum_40_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_18( .activation_in(reg_activation_40_17), .weight_in(reg_weight_39_18), .partial_sum_in(reg_psum_39_18), .reg_activation(reg_activation_40_18), .reg_weight(reg_weight_40_18), .reg_partial_sum(reg_psum_40_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_19( .activation_in(reg_activation_40_18), .weight_in(reg_weight_39_19), .partial_sum_in(reg_psum_39_19), .reg_activation(reg_activation_40_19), .reg_weight(reg_weight_40_19), .reg_partial_sum(reg_psum_40_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_20( .activation_in(reg_activation_40_19), .weight_in(reg_weight_39_20), .partial_sum_in(reg_psum_39_20), .reg_activation(reg_activation_40_20), .reg_weight(reg_weight_40_20), .reg_partial_sum(reg_psum_40_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_21( .activation_in(reg_activation_40_20), .weight_in(reg_weight_39_21), .partial_sum_in(reg_psum_39_21), .reg_activation(reg_activation_40_21), .reg_weight(reg_weight_40_21), .reg_partial_sum(reg_psum_40_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_22( .activation_in(reg_activation_40_21), .weight_in(reg_weight_39_22), .partial_sum_in(reg_psum_39_22), .reg_activation(reg_activation_40_22), .reg_weight(reg_weight_40_22), .reg_partial_sum(reg_psum_40_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_23( .activation_in(reg_activation_40_22), .weight_in(reg_weight_39_23), .partial_sum_in(reg_psum_39_23), .reg_activation(reg_activation_40_23), .reg_weight(reg_weight_40_23), .reg_partial_sum(reg_psum_40_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_24( .activation_in(reg_activation_40_23), .weight_in(reg_weight_39_24), .partial_sum_in(reg_psum_39_24), .reg_activation(reg_activation_40_24), .reg_weight(reg_weight_40_24), .reg_partial_sum(reg_psum_40_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_25( .activation_in(reg_activation_40_24), .weight_in(reg_weight_39_25), .partial_sum_in(reg_psum_39_25), .reg_activation(reg_activation_40_25), .reg_weight(reg_weight_40_25), .reg_partial_sum(reg_psum_40_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_26( .activation_in(reg_activation_40_25), .weight_in(reg_weight_39_26), .partial_sum_in(reg_psum_39_26), .reg_activation(reg_activation_40_26), .reg_weight(reg_weight_40_26), .reg_partial_sum(reg_psum_40_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_27( .activation_in(reg_activation_40_26), .weight_in(reg_weight_39_27), .partial_sum_in(reg_psum_39_27), .reg_activation(reg_activation_40_27), .reg_weight(reg_weight_40_27), .reg_partial_sum(reg_psum_40_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_28( .activation_in(reg_activation_40_27), .weight_in(reg_weight_39_28), .partial_sum_in(reg_psum_39_28), .reg_activation(reg_activation_40_28), .reg_weight(reg_weight_40_28), .reg_partial_sum(reg_psum_40_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_29( .activation_in(reg_activation_40_28), .weight_in(reg_weight_39_29), .partial_sum_in(reg_psum_39_29), .reg_activation(reg_activation_40_29), .reg_weight(reg_weight_40_29), .reg_partial_sum(reg_psum_40_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_30( .activation_in(reg_activation_40_29), .weight_in(reg_weight_39_30), .partial_sum_in(reg_psum_39_30), .reg_activation(reg_activation_40_30), .reg_weight(reg_weight_40_30), .reg_partial_sum(reg_psum_40_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_31( .activation_in(reg_activation_40_30), .weight_in(reg_weight_39_31), .partial_sum_in(reg_psum_39_31), .reg_activation(reg_activation_40_31), .reg_weight(reg_weight_40_31), .reg_partial_sum(reg_psum_40_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_32( .activation_in(reg_activation_40_31), .weight_in(reg_weight_39_32), .partial_sum_in(reg_psum_39_32), .reg_activation(reg_activation_40_32), .reg_weight(reg_weight_40_32), .reg_partial_sum(reg_psum_40_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_33( .activation_in(reg_activation_40_32), .weight_in(reg_weight_39_33), .partial_sum_in(reg_psum_39_33), .reg_activation(reg_activation_40_33), .reg_weight(reg_weight_40_33), .reg_partial_sum(reg_psum_40_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_34( .activation_in(reg_activation_40_33), .weight_in(reg_weight_39_34), .partial_sum_in(reg_psum_39_34), .reg_activation(reg_activation_40_34), .reg_weight(reg_weight_40_34), .reg_partial_sum(reg_psum_40_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_35( .activation_in(reg_activation_40_34), .weight_in(reg_weight_39_35), .partial_sum_in(reg_psum_39_35), .reg_activation(reg_activation_40_35), .reg_weight(reg_weight_40_35), .reg_partial_sum(reg_psum_40_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_36( .activation_in(reg_activation_40_35), .weight_in(reg_weight_39_36), .partial_sum_in(reg_psum_39_36), .reg_activation(reg_activation_40_36), .reg_weight(reg_weight_40_36), .reg_partial_sum(reg_psum_40_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_37( .activation_in(reg_activation_40_36), .weight_in(reg_weight_39_37), .partial_sum_in(reg_psum_39_37), .reg_activation(reg_activation_40_37), .reg_weight(reg_weight_40_37), .reg_partial_sum(reg_psum_40_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_38( .activation_in(reg_activation_40_37), .weight_in(reg_weight_39_38), .partial_sum_in(reg_psum_39_38), .reg_activation(reg_activation_40_38), .reg_weight(reg_weight_40_38), .reg_partial_sum(reg_psum_40_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_39( .activation_in(reg_activation_40_38), .weight_in(reg_weight_39_39), .partial_sum_in(reg_psum_39_39), .reg_activation(reg_activation_40_39), .reg_weight(reg_weight_40_39), .reg_partial_sum(reg_psum_40_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_40( .activation_in(reg_activation_40_39), .weight_in(reg_weight_39_40), .partial_sum_in(reg_psum_39_40), .reg_activation(reg_activation_40_40), .reg_weight(reg_weight_40_40), .reg_partial_sum(reg_psum_40_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_41( .activation_in(reg_activation_40_40), .weight_in(reg_weight_39_41), .partial_sum_in(reg_psum_39_41), .reg_activation(reg_activation_40_41), .reg_weight(reg_weight_40_41), .reg_partial_sum(reg_psum_40_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_42( .activation_in(reg_activation_40_41), .weight_in(reg_weight_39_42), .partial_sum_in(reg_psum_39_42), .reg_activation(reg_activation_40_42), .reg_weight(reg_weight_40_42), .reg_partial_sum(reg_psum_40_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_43( .activation_in(reg_activation_40_42), .weight_in(reg_weight_39_43), .partial_sum_in(reg_psum_39_43), .reg_activation(reg_activation_40_43), .reg_weight(reg_weight_40_43), .reg_partial_sum(reg_psum_40_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_44( .activation_in(reg_activation_40_43), .weight_in(reg_weight_39_44), .partial_sum_in(reg_psum_39_44), .reg_activation(reg_activation_40_44), .reg_weight(reg_weight_40_44), .reg_partial_sum(reg_psum_40_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_45( .activation_in(reg_activation_40_44), .weight_in(reg_weight_39_45), .partial_sum_in(reg_psum_39_45), .reg_activation(reg_activation_40_45), .reg_weight(reg_weight_40_45), .reg_partial_sum(reg_psum_40_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_46( .activation_in(reg_activation_40_45), .weight_in(reg_weight_39_46), .partial_sum_in(reg_psum_39_46), .reg_activation(reg_activation_40_46), .reg_weight(reg_weight_40_46), .reg_partial_sum(reg_psum_40_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_47( .activation_in(reg_activation_40_46), .weight_in(reg_weight_39_47), .partial_sum_in(reg_psum_39_47), .reg_activation(reg_activation_40_47), .reg_weight(reg_weight_40_47), .reg_partial_sum(reg_psum_40_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_48( .activation_in(reg_activation_40_47), .weight_in(reg_weight_39_48), .partial_sum_in(reg_psum_39_48), .reg_activation(reg_activation_40_48), .reg_weight(reg_weight_40_48), .reg_partial_sum(reg_psum_40_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_49( .activation_in(reg_activation_40_48), .weight_in(reg_weight_39_49), .partial_sum_in(reg_psum_39_49), .reg_activation(reg_activation_40_49), .reg_weight(reg_weight_40_49), .reg_partial_sum(reg_psum_40_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_50( .activation_in(reg_activation_40_49), .weight_in(reg_weight_39_50), .partial_sum_in(reg_psum_39_50), .reg_activation(reg_activation_40_50), .reg_weight(reg_weight_40_50), .reg_partial_sum(reg_psum_40_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_51( .activation_in(reg_activation_40_50), .weight_in(reg_weight_39_51), .partial_sum_in(reg_psum_39_51), .reg_activation(reg_activation_40_51), .reg_weight(reg_weight_40_51), .reg_partial_sum(reg_psum_40_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_52( .activation_in(reg_activation_40_51), .weight_in(reg_weight_39_52), .partial_sum_in(reg_psum_39_52), .reg_activation(reg_activation_40_52), .reg_weight(reg_weight_40_52), .reg_partial_sum(reg_psum_40_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_53( .activation_in(reg_activation_40_52), .weight_in(reg_weight_39_53), .partial_sum_in(reg_psum_39_53), .reg_activation(reg_activation_40_53), .reg_weight(reg_weight_40_53), .reg_partial_sum(reg_psum_40_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_54( .activation_in(reg_activation_40_53), .weight_in(reg_weight_39_54), .partial_sum_in(reg_psum_39_54), .reg_activation(reg_activation_40_54), .reg_weight(reg_weight_40_54), .reg_partial_sum(reg_psum_40_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_55( .activation_in(reg_activation_40_54), .weight_in(reg_weight_39_55), .partial_sum_in(reg_psum_39_55), .reg_activation(reg_activation_40_55), .reg_weight(reg_weight_40_55), .reg_partial_sum(reg_psum_40_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_56( .activation_in(reg_activation_40_55), .weight_in(reg_weight_39_56), .partial_sum_in(reg_psum_39_56), .reg_activation(reg_activation_40_56), .reg_weight(reg_weight_40_56), .reg_partial_sum(reg_psum_40_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_57( .activation_in(reg_activation_40_56), .weight_in(reg_weight_39_57), .partial_sum_in(reg_psum_39_57), .reg_activation(reg_activation_40_57), .reg_weight(reg_weight_40_57), .reg_partial_sum(reg_psum_40_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_58( .activation_in(reg_activation_40_57), .weight_in(reg_weight_39_58), .partial_sum_in(reg_psum_39_58), .reg_activation(reg_activation_40_58), .reg_weight(reg_weight_40_58), .reg_partial_sum(reg_psum_40_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_59( .activation_in(reg_activation_40_58), .weight_in(reg_weight_39_59), .partial_sum_in(reg_psum_39_59), .reg_activation(reg_activation_40_59), .reg_weight(reg_weight_40_59), .reg_partial_sum(reg_psum_40_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_60( .activation_in(reg_activation_40_59), .weight_in(reg_weight_39_60), .partial_sum_in(reg_psum_39_60), .reg_activation(reg_activation_40_60), .reg_weight(reg_weight_40_60), .reg_partial_sum(reg_psum_40_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_61( .activation_in(reg_activation_40_60), .weight_in(reg_weight_39_61), .partial_sum_in(reg_psum_39_61), .reg_activation(reg_activation_40_61), .reg_weight(reg_weight_40_61), .reg_partial_sum(reg_psum_40_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_62( .activation_in(reg_activation_40_61), .weight_in(reg_weight_39_62), .partial_sum_in(reg_psum_39_62), .reg_activation(reg_activation_40_62), .reg_weight(reg_weight_40_62), .reg_partial_sum(reg_psum_40_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U40_63( .activation_in(reg_activation_40_62), .weight_in(reg_weight_39_63), .partial_sum_in(reg_psum_39_63), .reg_weight(reg_weight_40_63), .reg_partial_sum(reg_psum_40_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_0( .activation_in(in_activation_41), .weight_in(reg_weight_40_0), .partial_sum_in(reg_psum_40_0), .reg_activation(reg_activation_41_0), .reg_weight(reg_weight_41_0), .reg_partial_sum(reg_psum_41_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_1( .activation_in(reg_activation_41_0), .weight_in(reg_weight_40_1), .partial_sum_in(reg_psum_40_1), .reg_activation(reg_activation_41_1), .reg_weight(reg_weight_41_1), .reg_partial_sum(reg_psum_41_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_2( .activation_in(reg_activation_41_1), .weight_in(reg_weight_40_2), .partial_sum_in(reg_psum_40_2), .reg_activation(reg_activation_41_2), .reg_weight(reg_weight_41_2), .reg_partial_sum(reg_psum_41_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_3( .activation_in(reg_activation_41_2), .weight_in(reg_weight_40_3), .partial_sum_in(reg_psum_40_3), .reg_activation(reg_activation_41_3), .reg_weight(reg_weight_41_3), .reg_partial_sum(reg_psum_41_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_4( .activation_in(reg_activation_41_3), .weight_in(reg_weight_40_4), .partial_sum_in(reg_psum_40_4), .reg_activation(reg_activation_41_4), .reg_weight(reg_weight_41_4), .reg_partial_sum(reg_psum_41_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_5( .activation_in(reg_activation_41_4), .weight_in(reg_weight_40_5), .partial_sum_in(reg_psum_40_5), .reg_activation(reg_activation_41_5), .reg_weight(reg_weight_41_5), .reg_partial_sum(reg_psum_41_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_6( .activation_in(reg_activation_41_5), .weight_in(reg_weight_40_6), .partial_sum_in(reg_psum_40_6), .reg_activation(reg_activation_41_6), .reg_weight(reg_weight_41_6), .reg_partial_sum(reg_psum_41_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_7( .activation_in(reg_activation_41_6), .weight_in(reg_weight_40_7), .partial_sum_in(reg_psum_40_7), .reg_activation(reg_activation_41_7), .reg_weight(reg_weight_41_7), .reg_partial_sum(reg_psum_41_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_8( .activation_in(reg_activation_41_7), .weight_in(reg_weight_40_8), .partial_sum_in(reg_psum_40_8), .reg_activation(reg_activation_41_8), .reg_weight(reg_weight_41_8), .reg_partial_sum(reg_psum_41_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_9( .activation_in(reg_activation_41_8), .weight_in(reg_weight_40_9), .partial_sum_in(reg_psum_40_9), .reg_activation(reg_activation_41_9), .reg_weight(reg_weight_41_9), .reg_partial_sum(reg_psum_41_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_10( .activation_in(reg_activation_41_9), .weight_in(reg_weight_40_10), .partial_sum_in(reg_psum_40_10), .reg_activation(reg_activation_41_10), .reg_weight(reg_weight_41_10), .reg_partial_sum(reg_psum_41_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_11( .activation_in(reg_activation_41_10), .weight_in(reg_weight_40_11), .partial_sum_in(reg_psum_40_11), .reg_activation(reg_activation_41_11), .reg_weight(reg_weight_41_11), .reg_partial_sum(reg_psum_41_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_12( .activation_in(reg_activation_41_11), .weight_in(reg_weight_40_12), .partial_sum_in(reg_psum_40_12), .reg_activation(reg_activation_41_12), .reg_weight(reg_weight_41_12), .reg_partial_sum(reg_psum_41_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_13( .activation_in(reg_activation_41_12), .weight_in(reg_weight_40_13), .partial_sum_in(reg_psum_40_13), .reg_activation(reg_activation_41_13), .reg_weight(reg_weight_41_13), .reg_partial_sum(reg_psum_41_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_14( .activation_in(reg_activation_41_13), .weight_in(reg_weight_40_14), .partial_sum_in(reg_psum_40_14), .reg_activation(reg_activation_41_14), .reg_weight(reg_weight_41_14), .reg_partial_sum(reg_psum_41_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_15( .activation_in(reg_activation_41_14), .weight_in(reg_weight_40_15), .partial_sum_in(reg_psum_40_15), .reg_activation(reg_activation_41_15), .reg_weight(reg_weight_41_15), .reg_partial_sum(reg_psum_41_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_16( .activation_in(reg_activation_41_15), .weight_in(reg_weight_40_16), .partial_sum_in(reg_psum_40_16), .reg_activation(reg_activation_41_16), .reg_weight(reg_weight_41_16), .reg_partial_sum(reg_psum_41_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_17( .activation_in(reg_activation_41_16), .weight_in(reg_weight_40_17), .partial_sum_in(reg_psum_40_17), .reg_activation(reg_activation_41_17), .reg_weight(reg_weight_41_17), .reg_partial_sum(reg_psum_41_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_18( .activation_in(reg_activation_41_17), .weight_in(reg_weight_40_18), .partial_sum_in(reg_psum_40_18), .reg_activation(reg_activation_41_18), .reg_weight(reg_weight_41_18), .reg_partial_sum(reg_psum_41_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_19( .activation_in(reg_activation_41_18), .weight_in(reg_weight_40_19), .partial_sum_in(reg_psum_40_19), .reg_activation(reg_activation_41_19), .reg_weight(reg_weight_41_19), .reg_partial_sum(reg_psum_41_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_20( .activation_in(reg_activation_41_19), .weight_in(reg_weight_40_20), .partial_sum_in(reg_psum_40_20), .reg_activation(reg_activation_41_20), .reg_weight(reg_weight_41_20), .reg_partial_sum(reg_psum_41_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_21( .activation_in(reg_activation_41_20), .weight_in(reg_weight_40_21), .partial_sum_in(reg_psum_40_21), .reg_activation(reg_activation_41_21), .reg_weight(reg_weight_41_21), .reg_partial_sum(reg_psum_41_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_22( .activation_in(reg_activation_41_21), .weight_in(reg_weight_40_22), .partial_sum_in(reg_psum_40_22), .reg_activation(reg_activation_41_22), .reg_weight(reg_weight_41_22), .reg_partial_sum(reg_psum_41_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_23( .activation_in(reg_activation_41_22), .weight_in(reg_weight_40_23), .partial_sum_in(reg_psum_40_23), .reg_activation(reg_activation_41_23), .reg_weight(reg_weight_41_23), .reg_partial_sum(reg_psum_41_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_24( .activation_in(reg_activation_41_23), .weight_in(reg_weight_40_24), .partial_sum_in(reg_psum_40_24), .reg_activation(reg_activation_41_24), .reg_weight(reg_weight_41_24), .reg_partial_sum(reg_psum_41_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_25( .activation_in(reg_activation_41_24), .weight_in(reg_weight_40_25), .partial_sum_in(reg_psum_40_25), .reg_activation(reg_activation_41_25), .reg_weight(reg_weight_41_25), .reg_partial_sum(reg_psum_41_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_26( .activation_in(reg_activation_41_25), .weight_in(reg_weight_40_26), .partial_sum_in(reg_psum_40_26), .reg_activation(reg_activation_41_26), .reg_weight(reg_weight_41_26), .reg_partial_sum(reg_psum_41_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_27( .activation_in(reg_activation_41_26), .weight_in(reg_weight_40_27), .partial_sum_in(reg_psum_40_27), .reg_activation(reg_activation_41_27), .reg_weight(reg_weight_41_27), .reg_partial_sum(reg_psum_41_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_28( .activation_in(reg_activation_41_27), .weight_in(reg_weight_40_28), .partial_sum_in(reg_psum_40_28), .reg_activation(reg_activation_41_28), .reg_weight(reg_weight_41_28), .reg_partial_sum(reg_psum_41_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_29( .activation_in(reg_activation_41_28), .weight_in(reg_weight_40_29), .partial_sum_in(reg_psum_40_29), .reg_activation(reg_activation_41_29), .reg_weight(reg_weight_41_29), .reg_partial_sum(reg_psum_41_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_30( .activation_in(reg_activation_41_29), .weight_in(reg_weight_40_30), .partial_sum_in(reg_psum_40_30), .reg_activation(reg_activation_41_30), .reg_weight(reg_weight_41_30), .reg_partial_sum(reg_psum_41_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_31( .activation_in(reg_activation_41_30), .weight_in(reg_weight_40_31), .partial_sum_in(reg_psum_40_31), .reg_activation(reg_activation_41_31), .reg_weight(reg_weight_41_31), .reg_partial_sum(reg_psum_41_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_32( .activation_in(reg_activation_41_31), .weight_in(reg_weight_40_32), .partial_sum_in(reg_psum_40_32), .reg_activation(reg_activation_41_32), .reg_weight(reg_weight_41_32), .reg_partial_sum(reg_psum_41_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_33( .activation_in(reg_activation_41_32), .weight_in(reg_weight_40_33), .partial_sum_in(reg_psum_40_33), .reg_activation(reg_activation_41_33), .reg_weight(reg_weight_41_33), .reg_partial_sum(reg_psum_41_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_34( .activation_in(reg_activation_41_33), .weight_in(reg_weight_40_34), .partial_sum_in(reg_psum_40_34), .reg_activation(reg_activation_41_34), .reg_weight(reg_weight_41_34), .reg_partial_sum(reg_psum_41_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_35( .activation_in(reg_activation_41_34), .weight_in(reg_weight_40_35), .partial_sum_in(reg_psum_40_35), .reg_activation(reg_activation_41_35), .reg_weight(reg_weight_41_35), .reg_partial_sum(reg_psum_41_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_36( .activation_in(reg_activation_41_35), .weight_in(reg_weight_40_36), .partial_sum_in(reg_psum_40_36), .reg_activation(reg_activation_41_36), .reg_weight(reg_weight_41_36), .reg_partial_sum(reg_psum_41_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_37( .activation_in(reg_activation_41_36), .weight_in(reg_weight_40_37), .partial_sum_in(reg_psum_40_37), .reg_activation(reg_activation_41_37), .reg_weight(reg_weight_41_37), .reg_partial_sum(reg_psum_41_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_38( .activation_in(reg_activation_41_37), .weight_in(reg_weight_40_38), .partial_sum_in(reg_psum_40_38), .reg_activation(reg_activation_41_38), .reg_weight(reg_weight_41_38), .reg_partial_sum(reg_psum_41_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_39( .activation_in(reg_activation_41_38), .weight_in(reg_weight_40_39), .partial_sum_in(reg_psum_40_39), .reg_activation(reg_activation_41_39), .reg_weight(reg_weight_41_39), .reg_partial_sum(reg_psum_41_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_40( .activation_in(reg_activation_41_39), .weight_in(reg_weight_40_40), .partial_sum_in(reg_psum_40_40), .reg_activation(reg_activation_41_40), .reg_weight(reg_weight_41_40), .reg_partial_sum(reg_psum_41_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_41( .activation_in(reg_activation_41_40), .weight_in(reg_weight_40_41), .partial_sum_in(reg_psum_40_41), .reg_activation(reg_activation_41_41), .reg_weight(reg_weight_41_41), .reg_partial_sum(reg_psum_41_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_42( .activation_in(reg_activation_41_41), .weight_in(reg_weight_40_42), .partial_sum_in(reg_psum_40_42), .reg_activation(reg_activation_41_42), .reg_weight(reg_weight_41_42), .reg_partial_sum(reg_psum_41_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_43( .activation_in(reg_activation_41_42), .weight_in(reg_weight_40_43), .partial_sum_in(reg_psum_40_43), .reg_activation(reg_activation_41_43), .reg_weight(reg_weight_41_43), .reg_partial_sum(reg_psum_41_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_44( .activation_in(reg_activation_41_43), .weight_in(reg_weight_40_44), .partial_sum_in(reg_psum_40_44), .reg_activation(reg_activation_41_44), .reg_weight(reg_weight_41_44), .reg_partial_sum(reg_psum_41_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_45( .activation_in(reg_activation_41_44), .weight_in(reg_weight_40_45), .partial_sum_in(reg_psum_40_45), .reg_activation(reg_activation_41_45), .reg_weight(reg_weight_41_45), .reg_partial_sum(reg_psum_41_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_46( .activation_in(reg_activation_41_45), .weight_in(reg_weight_40_46), .partial_sum_in(reg_psum_40_46), .reg_activation(reg_activation_41_46), .reg_weight(reg_weight_41_46), .reg_partial_sum(reg_psum_41_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_47( .activation_in(reg_activation_41_46), .weight_in(reg_weight_40_47), .partial_sum_in(reg_psum_40_47), .reg_activation(reg_activation_41_47), .reg_weight(reg_weight_41_47), .reg_partial_sum(reg_psum_41_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_48( .activation_in(reg_activation_41_47), .weight_in(reg_weight_40_48), .partial_sum_in(reg_psum_40_48), .reg_activation(reg_activation_41_48), .reg_weight(reg_weight_41_48), .reg_partial_sum(reg_psum_41_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_49( .activation_in(reg_activation_41_48), .weight_in(reg_weight_40_49), .partial_sum_in(reg_psum_40_49), .reg_activation(reg_activation_41_49), .reg_weight(reg_weight_41_49), .reg_partial_sum(reg_psum_41_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_50( .activation_in(reg_activation_41_49), .weight_in(reg_weight_40_50), .partial_sum_in(reg_psum_40_50), .reg_activation(reg_activation_41_50), .reg_weight(reg_weight_41_50), .reg_partial_sum(reg_psum_41_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_51( .activation_in(reg_activation_41_50), .weight_in(reg_weight_40_51), .partial_sum_in(reg_psum_40_51), .reg_activation(reg_activation_41_51), .reg_weight(reg_weight_41_51), .reg_partial_sum(reg_psum_41_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_52( .activation_in(reg_activation_41_51), .weight_in(reg_weight_40_52), .partial_sum_in(reg_psum_40_52), .reg_activation(reg_activation_41_52), .reg_weight(reg_weight_41_52), .reg_partial_sum(reg_psum_41_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_53( .activation_in(reg_activation_41_52), .weight_in(reg_weight_40_53), .partial_sum_in(reg_psum_40_53), .reg_activation(reg_activation_41_53), .reg_weight(reg_weight_41_53), .reg_partial_sum(reg_psum_41_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_54( .activation_in(reg_activation_41_53), .weight_in(reg_weight_40_54), .partial_sum_in(reg_psum_40_54), .reg_activation(reg_activation_41_54), .reg_weight(reg_weight_41_54), .reg_partial_sum(reg_psum_41_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_55( .activation_in(reg_activation_41_54), .weight_in(reg_weight_40_55), .partial_sum_in(reg_psum_40_55), .reg_activation(reg_activation_41_55), .reg_weight(reg_weight_41_55), .reg_partial_sum(reg_psum_41_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_56( .activation_in(reg_activation_41_55), .weight_in(reg_weight_40_56), .partial_sum_in(reg_psum_40_56), .reg_activation(reg_activation_41_56), .reg_weight(reg_weight_41_56), .reg_partial_sum(reg_psum_41_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_57( .activation_in(reg_activation_41_56), .weight_in(reg_weight_40_57), .partial_sum_in(reg_psum_40_57), .reg_activation(reg_activation_41_57), .reg_weight(reg_weight_41_57), .reg_partial_sum(reg_psum_41_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_58( .activation_in(reg_activation_41_57), .weight_in(reg_weight_40_58), .partial_sum_in(reg_psum_40_58), .reg_activation(reg_activation_41_58), .reg_weight(reg_weight_41_58), .reg_partial_sum(reg_psum_41_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_59( .activation_in(reg_activation_41_58), .weight_in(reg_weight_40_59), .partial_sum_in(reg_psum_40_59), .reg_activation(reg_activation_41_59), .reg_weight(reg_weight_41_59), .reg_partial_sum(reg_psum_41_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_60( .activation_in(reg_activation_41_59), .weight_in(reg_weight_40_60), .partial_sum_in(reg_psum_40_60), .reg_activation(reg_activation_41_60), .reg_weight(reg_weight_41_60), .reg_partial_sum(reg_psum_41_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_61( .activation_in(reg_activation_41_60), .weight_in(reg_weight_40_61), .partial_sum_in(reg_psum_40_61), .reg_activation(reg_activation_41_61), .reg_weight(reg_weight_41_61), .reg_partial_sum(reg_psum_41_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_62( .activation_in(reg_activation_41_61), .weight_in(reg_weight_40_62), .partial_sum_in(reg_psum_40_62), .reg_activation(reg_activation_41_62), .reg_weight(reg_weight_41_62), .reg_partial_sum(reg_psum_41_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U41_63( .activation_in(reg_activation_41_62), .weight_in(reg_weight_40_63), .partial_sum_in(reg_psum_40_63), .reg_weight(reg_weight_41_63), .reg_partial_sum(reg_psum_41_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_0( .activation_in(in_activation_42), .weight_in(reg_weight_41_0), .partial_sum_in(reg_psum_41_0), .reg_activation(reg_activation_42_0), .reg_weight(reg_weight_42_0), .reg_partial_sum(reg_psum_42_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_1( .activation_in(reg_activation_42_0), .weight_in(reg_weight_41_1), .partial_sum_in(reg_psum_41_1), .reg_activation(reg_activation_42_1), .reg_weight(reg_weight_42_1), .reg_partial_sum(reg_psum_42_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_2( .activation_in(reg_activation_42_1), .weight_in(reg_weight_41_2), .partial_sum_in(reg_psum_41_2), .reg_activation(reg_activation_42_2), .reg_weight(reg_weight_42_2), .reg_partial_sum(reg_psum_42_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_3( .activation_in(reg_activation_42_2), .weight_in(reg_weight_41_3), .partial_sum_in(reg_psum_41_3), .reg_activation(reg_activation_42_3), .reg_weight(reg_weight_42_3), .reg_partial_sum(reg_psum_42_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_4( .activation_in(reg_activation_42_3), .weight_in(reg_weight_41_4), .partial_sum_in(reg_psum_41_4), .reg_activation(reg_activation_42_4), .reg_weight(reg_weight_42_4), .reg_partial_sum(reg_psum_42_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_5( .activation_in(reg_activation_42_4), .weight_in(reg_weight_41_5), .partial_sum_in(reg_psum_41_5), .reg_activation(reg_activation_42_5), .reg_weight(reg_weight_42_5), .reg_partial_sum(reg_psum_42_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_6( .activation_in(reg_activation_42_5), .weight_in(reg_weight_41_6), .partial_sum_in(reg_psum_41_6), .reg_activation(reg_activation_42_6), .reg_weight(reg_weight_42_6), .reg_partial_sum(reg_psum_42_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_7( .activation_in(reg_activation_42_6), .weight_in(reg_weight_41_7), .partial_sum_in(reg_psum_41_7), .reg_activation(reg_activation_42_7), .reg_weight(reg_weight_42_7), .reg_partial_sum(reg_psum_42_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_8( .activation_in(reg_activation_42_7), .weight_in(reg_weight_41_8), .partial_sum_in(reg_psum_41_8), .reg_activation(reg_activation_42_8), .reg_weight(reg_weight_42_8), .reg_partial_sum(reg_psum_42_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_9( .activation_in(reg_activation_42_8), .weight_in(reg_weight_41_9), .partial_sum_in(reg_psum_41_9), .reg_activation(reg_activation_42_9), .reg_weight(reg_weight_42_9), .reg_partial_sum(reg_psum_42_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_10( .activation_in(reg_activation_42_9), .weight_in(reg_weight_41_10), .partial_sum_in(reg_psum_41_10), .reg_activation(reg_activation_42_10), .reg_weight(reg_weight_42_10), .reg_partial_sum(reg_psum_42_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_11( .activation_in(reg_activation_42_10), .weight_in(reg_weight_41_11), .partial_sum_in(reg_psum_41_11), .reg_activation(reg_activation_42_11), .reg_weight(reg_weight_42_11), .reg_partial_sum(reg_psum_42_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_12( .activation_in(reg_activation_42_11), .weight_in(reg_weight_41_12), .partial_sum_in(reg_psum_41_12), .reg_activation(reg_activation_42_12), .reg_weight(reg_weight_42_12), .reg_partial_sum(reg_psum_42_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_13( .activation_in(reg_activation_42_12), .weight_in(reg_weight_41_13), .partial_sum_in(reg_psum_41_13), .reg_activation(reg_activation_42_13), .reg_weight(reg_weight_42_13), .reg_partial_sum(reg_psum_42_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_14( .activation_in(reg_activation_42_13), .weight_in(reg_weight_41_14), .partial_sum_in(reg_psum_41_14), .reg_activation(reg_activation_42_14), .reg_weight(reg_weight_42_14), .reg_partial_sum(reg_psum_42_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_15( .activation_in(reg_activation_42_14), .weight_in(reg_weight_41_15), .partial_sum_in(reg_psum_41_15), .reg_activation(reg_activation_42_15), .reg_weight(reg_weight_42_15), .reg_partial_sum(reg_psum_42_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_16( .activation_in(reg_activation_42_15), .weight_in(reg_weight_41_16), .partial_sum_in(reg_psum_41_16), .reg_activation(reg_activation_42_16), .reg_weight(reg_weight_42_16), .reg_partial_sum(reg_psum_42_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_17( .activation_in(reg_activation_42_16), .weight_in(reg_weight_41_17), .partial_sum_in(reg_psum_41_17), .reg_activation(reg_activation_42_17), .reg_weight(reg_weight_42_17), .reg_partial_sum(reg_psum_42_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_18( .activation_in(reg_activation_42_17), .weight_in(reg_weight_41_18), .partial_sum_in(reg_psum_41_18), .reg_activation(reg_activation_42_18), .reg_weight(reg_weight_42_18), .reg_partial_sum(reg_psum_42_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_19( .activation_in(reg_activation_42_18), .weight_in(reg_weight_41_19), .partial_sum_in(reg_psum_41_19), .reg_activation(reg_activation_42_19), .reg_weight(reg_weight_42_19), .reg_partial_sum(reg_psum_42_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_20( .activation_in(reg_activation_42_19), .weight_in(reg_weight_41_20), .partial_sum_in(reg_psum_41_20), .reg_activation(reg_activation_42_20), .reg_weight(reg_weight_42_20), .reg_partial_sum(reg_psum_42_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_21( .activation_in(reg_activation_42_20), .weight_in(reg_weight_41_21), .partial_sum_in(reg_psum_41_21), .reg_activation(reg_activation_42_21), .reg_weight(reg_weight_42_21), .reg_partial_sum(reg_psum_42_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_22( .activation_in(reg_activation_42_21), .weight_in(reg_weight_41_22), .partial_sum_in(reg_psum_41_22), .reg_activation(reg_activation_42_22), .reg_weight(reg_weight_42_22), .reg_partial_sum(reg_psum_42_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_23( .activation_in(reg_activation_42_22), .weight_in(reg_weight_41_23), .partial_sum_in(reg_psum_41_23), .reg_activation(reg_activation_42_23), .reg_weight(reg_weight_42_23), .reg_partial_sum(reg_psum_42_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_24( .activation_in(reg_activation_42_23), .weight_in(reg_weight_41_24), .partial_sum_in(reg_psum_41_24), .reg_activation(reg_activation_42_24), .reg_weight(reg_weight_42_24), .reg_partial_sum(reg_psum_42_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_25( .activation_in(reg_activation_42_24), .weight_in(reg_weight_41_25), .partial_sum_in(reg_psum_41_25), .reg_activation(reg_activation_42_25), .reg_weight(reg_weight_42_25), .reg_partial_sum(reg_psum_42_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_26( .activation_in(reg_activation_42_25), .weight_in(reg_weight_41_26), .partial_sum_in(reg_psum_41_26), .reg_activation(reg_activation_42_26), .reg_weight(reg_weight_42_26), .reg_partial_sum(reg_psum_42_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_27( .activation_in(reg_activation_42_26), .weight_in(reg_weight_41_27), .partial_sum_in(reg_psum_41_27), .reg_activation(reg_activation_42_27), .reg_weight(reg_weight_42_27), .reg_partial_sum(reg_psum_42_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_28( .activation_in(reg_activation_42_27), .weight_in(reg_weight_41_28), .partial_sum_in(reg_psum_41_28), .reg_activation(reg_activation_42_28), .reg_weight(reg_weight_42_28), .reg_partial_sum(reg_psum_42_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_29( .activation_in(reg_activation_42_28), .weight_in(reg_weight_41_29), .partial_sum_in(reg_psum_41_29), .reg_activation(reg_activation_42_29), .reg_weight(reg_weight_42_29), .reg_partial_sum(reg_psum_42_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_30( .activation_in(reg_activation_42_29), .weight_in(reg_weight_41_30), .partial_sum_in(reg_psum_41_30), .reg_activation(reg_activation_42_30), .reg_weight(reg_weight_42_30), .reg_partial_sum(reg_psum_42_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_31( .activation_in(reg_activation_42_30), .weight_in(reg_weight_41_31), .partial_sum_in(reg_psum_41_31), .reg_activation(reg_activation_42_31), .reg_weight(reg_weight_42_31), .reg_partial_sum(reg_psum_42_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_32( .activation_in(reg_activation_42_31), .weight_in(reg_weight_41_32), .partial_sum_in(reg_psum_41_32), .reg_activation(reg_activation_42_32), .reg_weight(reg_weight_42_32), .reg_partial_sum(reg_psum_42_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_33( .activation_in(reg_activation_42_32), .weight_in(reg_weight_41_33), .partial_sum_in(reg_psum_41_33), .reg_activation(reg_activation_42_33), .reg_weight(reg_weight_42_33), .reg_partial_sum(reg_psum_42_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_34( .activation_in(reg_activation_42_33), .weight_in(reg_weight_41_34), .partial_sum_in(reg_psum_41_34), .reg_activation(reg_activation_42_34), .reg_weight(reg_weight_42_34), .reg_partial_sum(reg_psum_42_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_35( .activation_in(reg_activation_42_34), .weight_in(reg_weight_41_35), .partial_sum_in(reg_psum_41_35), .reg_activation(reg_activation_42_35), .reg_weight(reg_weight_42_35), .reg_partial_sum(reg_psum_42_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_36( .activation_in(reg_activation_42_35), .weight_in(reg_weight_41_36), .partial_sum_in(reg_psum_41_36), .reg_activation(reg_activation_42_36), .reg_weight(reg_weight_42_36), .reg_partial_sum(reg_psum_42_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_37( .activation_in(reg_activation_42_36), .weight_in(reg_weight_41_37), .partial_sum_in(reg_psum_41_37), .reg_activation(reg_activation_42_37), .reg_weight(reg_weight_42_37), .reg_partial_sum(reg_psum_42_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_38( .activation_in(reg_activation_42_37), .weight_in(reg_weight_41_38), .partial_sum_in(reg_psum_41_38), .reg_activation(reg_activation_42_38), .reg_weight(reg_weight_42_38), .reg_partial_sum(reg_psum_42_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_39( .activation_in(reg_activation_42_38), .weight_in(reg_weight_41_39), .partial_sum_in(reg_psum_41_39), .reg_activation(reg_activation_42_39), .reg_weight(reg_weight_42_39), .reg_partial_sum(reg_psum_42_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_40( .activation_in(reg_activation_42_39), .weight_in(reg_weight_41_40), .partial_sum_in(reg_psum_41_40), .reg_activation(reg_activation_42_40), .reg_weight(reg_weight_42_40), .reg_partial_sum(reg_psum_42_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_41( .activation_in(reg_activation_42_40), .weight_in(reg_weight_41_41), .partial_sum_in(reg_psum_41_41), .reg_activation(reg_activation_42_41), .reg_weight(reg_weight_42_41), .reg_partial_sum(reg_psum_42_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_42( .activation_in(reg_activation_42_41), .weight_in(reg_weight_41_42), .partial_sum_in(reg_psum_41_42), .reg_activation(reg_activation_42_42), .reg_weight(reg_weight_42_42), .reg_partial_sum(reg_psum_42_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_43( .activation_in(reg_activation_42_42), .weight_in(reg_weight_41_43), .partial_sum_in(reg_psum_41_43), .reg_activation(reg_activation_42_43), .reg_weight(reg_weight_42_43), .reg_partial_sum(reg_psum_42_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_44( .activation_in(reg_activation_42_43), .weight_in(reg_weight_41_44), .partial_sum_in(reg_psum_41_44), .reg_activation(reg_activation_42_44), .reg_weight(reg_weight_42_44), .reg_partial_sum(reg_psum_42_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_45( .activation_in(reg_activation_42_44), .weight_in(reg_weight_41_45), .partial_sum_in(reg_psum_41_45), .reg_activation(reg_activation_42_45), .reg_weight(reg_weight_42_45), .reg_partial_sum(reg_psum_42_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_46( .activation_in(reg_activation_42_45), .weight_in(reg_weight_41_46), .partial_sum_in(reg_psum_41_46), .reg_activation(reg_activation_42_46), .reg_weight(reg_weight_42_46), .reg_partial_sum(reg_psum_42_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_47( .activation_in(reg_activation_42_46), .weight_in(reg_weight_41_47), .partial_sum_in(reg_psum_41_47), .reg_activation(reg_activation_42_47), .reg_weight(reg_weight_42_47), .reg_partial_sum(reg_psum_42_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_48( .activation_in(reg_activation_42_47), .weight_in(reg_weight_41_48), .partial_sum_in(reg_psum_41_48), .reg_activation(reg_activation_42_48), .reg_weight(reg_weight_42_48), .reg_partial_sum(reg_psum_42_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_49( .activation_in(reg_activation_42_48), .weight_in(reg_weight_41_49), .partial_sum_in(reg_psum_41_49), .reg_activation(reg_activation_42_49), .reg_weight(reg_weight_42_49), .reg_partial_sum(reg_psum_42_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_50( .activation_in(reg_activation_42_49), .weight_in(reg_weight_41_50), .partial_sum_in(reg_psum_41_50), .reg_activation(reg_activation_42_50), .reg_weight(reg_weight_42_50), .reg_partial_sum(reg_psum_42_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_51( .activation_in(reg_activation_42_50), .weight_in(reg_weight_41_51), .partial_sum_in(reg_psum_41_51), .reg_activation(reg_activation_42_51), .reg_weight(reg_weight_42_51), .reg_partial_sum(reg_psum_42_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_52( .activation_in(reg_activation_42_51), .weight_in(reg_weight_41_52), .partial_sum_in(reg_psum_41_52), .reg_activation(reg_activation_42_52), .reg_weight(reg_weight_42_52), .reg_partial_sum(reg_psum_42_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_53( .activation_in(reg_activation_42_52), .weight_in(reg_weight_41_53), .partial_sum_in(reg_psum_41_53), .reg_activation(reg_activation_42_53), .reg_weight(reg_weight_42_53), .reg_partial_sum(reg_psum_42_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_54( .activation_in(reg_activation_42_53), .weight_in(reg_weight_41_54), .partial_sum_in(reg_psum_41_54), .reg_activation(reg_activation_42_54), .reg_weight(reg_weight_42_54), .reg_partial_sum(reg_psum_42_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_55( .activation_in(reg_activation_42_54), .weight_in(reg_weight_41_55), .partial_sum_in(reg_psum_41_55), .reg_activation(reg_activation_42_55), .reg_weight(reg_weight_42_55), .reg_partial_sum(reg_psum_42_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_56( .activation_in(reg_activation_42_55), .weight_in(reg_weight_41_56), .partial_sum_in(reg_psum_41_56), .reg_activation(reg_activation_42_56), .reg_weight(reg_weight_42_56), .reg_partial_sum(reg_psum_42_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_57( .activation_in(reg_activation_42_56), .weight_in(reg_weight_41_57), .partial_sum_in(reg_psum_41_57), .reg_activation(reg_activation_42_57), .reg_weight(reg_weight_42_57), .reg_partial_sum(reg_psum_42_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_58( .activation_in(reg_activation_42_57), .weight_in(reg_weight_41_58), .partial_sum_in(reg_psum_41_58), .reg_activation(reg_activation_42_58), .reg_weight(reg_weight_42_58), .reg_partial_sum(reg_psum_42_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_59( .activation_in(reg_activation_42_58), .weight_in(reg_weight_41_59), .partial_sum_in(reg_psum_41_59), .reg_activation(reg_activation_42_59), .reg_weight(reg_weight_42_59), .reg_partial_sum(reg_psum_42_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_60( .activation_in(reg_activation_42_59), .weight_in(reg_weight_41_60), .partial_sum_in(reg_psum_41_60), .reg_activation(reg_activation_42_60), .reg_weight(reg_weight_42_60), .reg_partial_sum(reg_psum_42_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_61( .activation_in(reg_activation_42_60), .weight_in(reg_weight_41_61), .partial_sum_in(reg_psum_41_61), .reg_activation(reg_activation_42_61), .reg_weight(reg_weight_42_61), .reg_partial_sum(reg_psum_42_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_62( .activation_in(reg_activation_42_61), .weight_in(reg_weight_41_62), .partial_sum_in(reg_psum_41_62), .reg_activation(reg_activation_42_62), .reg_weight(reg_weight_42_62), .reg_partial_sum(reg_psum_42_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U42_63( .activation_in(reg_activation_42_62), .weight_in(reg_weight_41_63), .partial_sum_in(reg_psum_41_63), .reg_weight(reg_weight_42_63), .reg_partial_sum(reg_psum_42_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_0( .activation_in(in_activation_43), .weight_in(reg_weight_42_0), .partial_sum_in(reg_psum_42_0), .reg_activation(reg_activation_43_0), .reg_weight(reg_weight_43_0), .reg_partial_sum(reg_psum_43_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_1( .activation_in(reg_activation_43_0), .weight_in(reg_weight_42_1), .partial_sum_in(reg_psum_42_1), .reg_activation(reg_activation_43_1), .reg_weight(reg_weight_43_1), .reg_partial_sum(reg_psum_43_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_2( .activation_in(reg_activation_43_1), .weight_in(reg_weight_42_2), .partial_sum_in(reg_psum_42_2), .reg_activation(reg_activation_43_2), .reg_weight(reg_weight_43_2), .reg_partial_sum(reg_psum_43_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_3( .activation_in(reg_activation_43_2), .weight_in(reg_weight_42_3), .partial_sum_in(reg_psum_42_3), .reg_activation(reg_activation_43_3), .reg_weight(reg_weight_43_3), .reg_partial_sum(reg_psum_43_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_4( .activation_in(reg_activation_43_3), .weight_in(reg_weight_42_4), .partial_sum_in(reg_psum_42_4), .reg_activation(reg_activation_43_4), .reg_weight(reg_weight_43_4), .reg_partial_sum(reg_psum_43_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_5( .activation_in(reg_activation_43_4), .weight_in(reg_weight_42_5), .partial_sum_in(reg_psum_42_5), .reg_activation(reg_activation_43_5), .reg_weight(reg_weight_43_5), .reg_partial_sum(reg_psum_43_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_6( .activation_in(reg_activation_43_5), .weight_in(reg_weight_42_6), .partial_sum_in(reg_psum_42_6), .reg_activation(reg_activation_43_6), .reg_weight(reg_weight_43_6), .reg_partial_sum(reg_psum_43_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_7( .activation_in(reg_activation_43_6), .weight_in(reg_weight_42_7), .partial_sum_in(reg_psum_42_7), .reg_activation(reg_activation_43_7), .reg_weight(reg_weight_43_7), .reg_partial_sum(reg_psum_43_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_8( .activation_in(reg_activation_43_7), .weight_in(reg_weight_42_8), .partial_sum_in(reg_psum_42_8), .reg_activation(reg_activation_43_8), .reg_weight(reg_weight_43_8), .reg_partial_sum(reg_psum_43_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_9( .activation_in(reg_activation_43_8), .weight_in(reg_weight_42_9), .partial_sum_in(reg_psum_42_9), .reg_activation(reg_activation_43_9), .reg_weight(reg_weight_43_9), .reg_partial_sum(reg_psum_43_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_10( .activation_in(reg_activation_43_9), .weight_in(reg_weight_42_10), .partial_sum_in(reg_psum_42_10), .reg_activation(reg_activation_43_10), .reg_weight(reg_weight_43_10), .reg_partial_sum(reg_psum_43_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_11( .activation_in(reg_activation_43_10), .weight_in(reg_weight_42_11), .partial_sum_in(reg_psum_42_11), .reg_activation(reg_activation_43_11), .reg_weight(reg_weight_43_11), .reg_partial_sum(reg_psum_43_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_12( .activation_in(reg_activation_43_11), .weight_in(reg_weight_42_12), .partial_sum_in(reg_psum_42_12), .reg_activation(reg_activation_43_12), .reg_weight(reg_weight_43_12), .reg_partial_sum(reg_psum_43_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_13( .activation_in(reg_activation_43_12), .weight_in(reg_weight_42_13), .partial_sum_in(reg_psum_42_13), .reg_activation(reg_activation_43_13), .reg_weight(reg_weight_43_13), .reg_partial_sum(reg_psum_43_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_14( .activation_in(reg_activation_43_13), .weight_in(reg_weight_42_14), .partial_sum_in(reg_psum_42_14), .reg_activation(reg_activation_43_14), .reg_weight(reg_weight_43_14), .reg_partial_sum(reg_psum_43_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_15( .activation_in(reg_activation_43_14), .weight_in(reg_weight_42_15), .partial_sum_in(reg_psum_42_15), .reg_activation(reg_activation_43_15), .reg_weight(reg_weight_43_15), .reg_partial_sum(reg_psum_43_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_16( .activation_in(reg_activation_43_15), .weight_in(reg_weight_42_16), .partial_sum_in(reg_psum_42_16), .reg_activation(reg_activation_43_16), .reg_weight(reg_weight_43_16), .reg_partial_sum(reg_psum_43_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_17( .activation_in(reg_activation_43_16), .weight_in(reg_weight_42_17), .partial_sum_in(reg_psum_42_17), .reg_activation(reg_activation_43_17), .reg_weight(reg_weight_43_17), .reg_partial_sum(reg_psum_43_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_18( .activation_in(reg_activation_43_17), .weight_in(reg_weight_42_18), .partial_sum_in(reg_psum_42_18), .reg_activation(reg_activation_43_18), .reg_weight(reg_weight_43_18), .reg_partial_sum(reg_psum_43_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_19( .activation_in(reg_activation_43_18), .weight_in(reg_weight_42_19), .partial_sum_in(reg_psum_42_19), .reg_activation(reg_activation_43_19), .reg_weight(reg_weight_43_19), .reg_partial_sum(reg_psum_43_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_20( .activation_in(reg_activation_43_19), .weight_in(reg_weight_42_20), .partial_sum_in(reg_psum_42_20), .reg_activation(reg_activation_43_20), .reg_weight(reg_weight_43_20), .reg_partial_sum(reg_psum_43_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_21( .activation_in(reg_activation_43_20), .weight_in(reg_weight_42_21), .partial_sum_in(reg_psum_42_21), .reg_activation(reg_activation_43_21), .reg_weight(reg_weight_43_21), .reg_partial_sum(reg_psum_43_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_22( .activation_in(reg_activation_43_21), .weight_in(reg_weight_42_22), .partial_sum_in(reg_psum_42_22), .reg_activation(reg_activation_43_22), .reg_weight(reg_weight_43_22), .reg_partial_sum(reg_psum_43_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_23( .activation_in(reg_activation_43_22), .weight_in(reg_weight_42_23), .partial_sum_in(reg_psum_42_23), .reg_activation(reg_activation_43_23), .reg_weight(reg_weight_43_23), .reg_partial_sum(reg_psum_43_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_24( .activation_in(reg_activation_43_23), .weight_in(reg_weight_42_24), .partial_sum_in(reg_psum_42_24), .reg_activation(reg_activation_43_24), .reg_weight(reg_weight_43_24), .reg_partial_sum(reg_psum_43_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_25( .activation_in(reg_activation_43_24), .weight_in(reg_weight_42_25), .partial_sum_in(reg_psum_42_25), .reg_activation(reg_activation_43_25), .reg_weight(reg_weight_43_25), .reg_partial_sum(reg_psum_43_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_26( .activation_in(reg_activation_43_25), .weight_in(reg_weight_42_26), .partial_sum_in(reg_psum_42_26), .reg_activation(reg_activation_43_26), .reg_weight(reg_weight_43_26), .reg_partial_sum(reg_psum_43_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_27( .activation_in(reg_activation_43_26), .weight_in(reg_weight_42_27), .partial_sum_in(reg_psum_42_27), .reg_activation(reg_activation_43_27), .reg_weight(reg_weight_43_27), .reg_partial_sum(reg_psum_43_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_28( .activation_in(reg_activation_43_27), .weight_in(reg_weight_42_28), .partial_sum_in(reg_psum_42_28), .reg_activation(reg_activation_43_28), .reg_weight(reg_weight_43_28), .reg_partial_sum(reg_psum_43_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_29( .activation_in(reg_activation_43_28), .weight_in(reg_weight_42_29), .partial_sum_in(reg_psum_42_29), .reg_activation(reg_activation_43_29), .reg_weight(reg_weight_43_29), .reg_partial_sum(reg_psum_43_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_30( .activation_in(reg_activation_43_29), .weight_in(reg_weight_42_30), .partial_sum_in(reg_psum_42_30), .reg_activation(reg_activation_43_30), .reg_weight(reg_weight_43_30), .reg_partial_sum(reg_psum_43_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_31( .activation_in(reg_activation_43_30), .weight_in(reg_weight_42_31), .partial_sum_in(reg_psum_42_31), .reg_activation(reg_activation_43_31), .reg_weight(reg_weight_43_31), .reg_partial_sum(reg_psum_43_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_32( .activation_in(reg_activation_43_31), .weight_in(reg_weight_42_32), .partial_sum_in(reg_psum_42_32), .reg_activation(reg_activation_43_32), .reg_weight(reg_weight_43_32), .reg_partial_sum(reg_psum_43_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_33( .activation_in(reg_activation_43_32), .weight_in(reg_weight_42_33), .partial_sum_in(reg_psum_42_33), .reg_activation(reg_activation_43_33), .reg_weight(reg_weight_43_33), .reg_partial_sum(reg_psum_43_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_34( .activation_in(reg_activation_43_33), .weight_in(reg_weight_42_34), .partial_sum_in(reg_psum_42_34), .reg_activation(reg_activation_43_34), .reg_weight(reg_weight_43_34), .reg_partial_sum(reg_psum_43_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_35( .activation_in(reg_activation_43_34), .weight_in(reg_weight_42_35), .partial_sum_in(reg_psum_42_35), .reg_activation(reg_activation_43_35), .reg_weight(reg_weight_43_35), .reg_partial_sum(reg_psum_43_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_36( .activation_in(reg_activation_43_35), .weight_in(reg_weight_42_36), .partial_sum_in(reg_psum_42_36), .reg_activation(reg_activation_43_36), .reg_weight(reg_weight_43_36), .reg_partial_sum(reg_psum_43_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_37( .activation_in(reg_activation_43_36), .weight_in(reg_weight_42_37), .partial_sum_in(reg_psum_42_37), .reg_activation(reg_activation_43_37), .reg_weight(reg_weight_43_37), .reg_partial_sum(reg_psum_43_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_38( .activation_in(reg_activation_43_37), .weight_in(reg_weight_42_38), .partial_sum_in(reg_psum_42_38), .reg_activation(reg_activation_43_38), .reg_weight(reg_weight_43_38), .reg_partial_sum(reg_psum_43_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_39( .activation_in(reg_activation_43_38), .weight_in(reg_weight_42_39), .partial_sum_in(reg_psum_42_39), .reg_activation(reg_activation_43_39), .reg_weight(reg_weight_43_39), .reg_partial_sum(reg_psum_43_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_40( .activation_in(reg_activation_43_39), .weight_in(reg_weight_42_40), .partial_sum_in(reg_psum_42_40), .reg_activation(reg_activation_43_40), .reg_weight(reg_weight_43_40), .reg_partial_sum(reg_psum_43_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_41( .activation_in(reg_activation_43_40), .weight_in(reg_weight_42_41), .partial_sum_in(reg_psum_42_41), .reg_activation(reg_activation_43_41), .reg_weight(reg_weight_43_41), .reg_partial_sum(reg_psum_43_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_42( .activation_in(reg_activation_43_41), .weight_in(reg_weight_42_42), .partial_sum_in(reg_psum_42_42), .reg_activation(reg_activation_43_42), .reg_weight(reg_weight_43_42), .reg_partial_sum(reg_psum_43_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_43( .activation_in(reg_activation_43_42), .weight_in(reg_weight_42_43), .partial_sum_in(reg_psum_42_43), .reg_activation(reg_activation_43_43), .reg_weight(reg_weight_43_43), .reg_partial_sum(reg_psum_43_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_44( .activation_in(reg_activation_43_43), .weight_in(reg_weight_42_44), .partial_sum_in(reg_psum_42_44), .reg_activation(reg_activation_43_44), .reg_weight(reg_weight_43_44), .reg_partial_sum(reg_psum_43_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_45( .activation_in(reg_activation_43_44), .weight_in(reg_weight_42_45), .partial_sum_in(reg_psum_42_45), .reg_activation(reg_activation_43_45), .reg_weight(reg_weight_43_45), .reg_partial_sum(reg_psum_43_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_46( .activation_in(reg_activation_43_45), .weight_in(reg_weight_42_46), .partial_sum_in(reg_psum_42_46), .reg_activation(reg_activation_43_46), .reg_weight(reg_weight_43_46), .reg_partial_sum(reg_psum_43_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_47( .activation_in(reg_activation_43_46), .weight_in(reg_weight_42_47), .partial_sum_in(reg_psum_42_47), .reg_activation(reg_activation_43_47), .reg_weight(reg_weight_43_47), .reg_partial_sum(reg_psum_43_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_48( .activation_in(reg_activation_43_47), .weight_in(reg_weight_42_48), .partial_sum_in(reg_psum_42_48), .reg_activation(reg_activation_43_48), .reg_weight(reg_weight_43_48), .reg_partial_sum(reg_psum_43_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_49( .activation_in(reg_activation_43_48), .weight_in(reg_weight_42_49), .partial_sum_in(reg_psum_42_49), .reg_activation(reg_activation_43_49), .reg_weight(reg_weight_43_49), .reg_partial_sum(reg_psum_43_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_50( .activation_in(reg_activation_43_49), .weight_in(reg_weight_42_50), .partial_sum_in(reg_psum_42_50), .reg_activation(reg_activation_43_50), .reg_weight(reg_weight_43_50), .reg_partial_sum(reg_psum_43_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_51( .activation_in(reg_activation_43_50), .weight_in(reg_weight_42_51), .partial_sum_in(reg_psum_42_51), .reg_activation(reg_activation_43_51), .reg_weight(reg_weight_43_51), .reg_partial_sum(reg_psum_43_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_52( .activation_in(reg_activation_43_51), .weight_in(reg_weight_42_52), .partial_sum_in(reg_psum_42_52), .reg_activation(reg_activation_43_52), .reg_weight(reg_weight_43_52), .reg_partial_sum(reg_psum_43_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_53( .activation_in(reg_activation_43_52), .weight_in(reg_weight_42_53), .partial_sum_in(reg_psum_42_53), .reg_activation(reg_activation_43_53), .reg_weight(reg_weight_43_53), .reg_partial_sum(reg_psum_43_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_54( .activation_in(reg_activation_43_53), .weight_in(reg_weight_42_54), .partial_sum_in(reg_psum_42_54), .reg_activation(reg_activation_43_54), .reg_weight(reg_weight_43_54), .reg_partial_sum(reg_psum_43_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_55( .activation_in(reg_activation_43_54), .weight_in(reg_weight_42_55), .partial_sum_in(reg_psum_42_55), .reg_activation(reg_activation_43_55), .reg_weight(reg_weight_43_55), .reg_partial_sum(reg_psum_43_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_56( .activation_in(reg_activation_43_55), .weight_in(reg_weight_42_56), .partial_sum_in(reg_psum_42_56), .reg_activation(reg_activation_43_56), .reg_weight(reg_weight_43_56), .reg_partial_sum(reg_psum_43_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_57( .activation_in(reg_activation_43_56), .weight_in(reg_weight_42_57), .partial_sum_in(reg_psum_42_57), .reg_activation(reg_activation_43_57), .reg_weight(reg_weight_43_57), .reg_partial_sum(reg_psum_43_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_58( .activation_in(reg_activation_43_57), .weight_in(reg_weight_42_58), .partial_sum_in(reg_psum_42_58), .reg_activation(reg_activation_43_58), .reg_weight(reg_weight_43_58), .reg_partial_sum(reg_psum_43_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_59( .activation_in(reg_activation_43_58), .weight_in(reg_weight_42_59), .partial_sum_in(reg_psum_42_59), .reg_activation(reg_activation_43_59), .reg_weight(reg_weight_43_59), .reg_partial_sum(reg_psum_43_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_60( .activation_in(reg_activation_43_59), .weight_in(reg_weight_42_60), .partial_sum_in(reg_psum_42_60), .reg_activation(reg_activation_43_60), .reg_weight(reg_weight_43_60), .reg_partial_sum(reg_psum_43_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_61( .activation_in(reg_activation_43_60), .weight_in(reg_weight_42_61), .partial_sum_in(reg_psum_42_61), .reg_activation(reg_activation_43_61), .reg_weight(reg_weight_43_61), .reg_partial_sum(reg_psum_43_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_62( .activation_in(reg_activation_43_61), .weight_in(reg_weight_42_62), .partial_sum_in(reg_psum_42_62), .reg_activation(reg_activation_43_62), .reg_weight(reg_weight_43_62), .reg_partial_sum(reg_psum_43_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U43_63( .activation_in(reg_activation_43_62), .weight_in(reg_weight_42_63), .partial_sum_in(reg_psum_42_63), .reg_weight(reg_weight_43_63), .reg_partial_sum(reg_psum_43_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_0( .activation_in(in_activation_44), .weight_in(reg_weight_43_0), .partial_sum_in(reg_psum_43_0), .reg_activation(reg_activation_44_0), .reg_weight(reg_weight_44_0), .reg_partial_sum(reg_psum_44_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_1( .activation_in(reg_activation_44_0), .weight_in(reg_weight_43_1), .partial_sum_in(reg_psum_43_1), .reg_activation(reg_activation_44_1), .reg_weight(reg_weight_44_1), .reg_partial_sum(reg_psum_44_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_2( .activation_in(reg_activation_44_1), .weight_in(reg_weight_43_2), .partial_sum_in(reg_psum_43_2), .reg_activation(reg_activation_44_2), .reg_weight(reg_weight_44_2), .reg_partial_sum(reg_psum_44_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_3( .activation_in(reg_activation_44_2), .weight_in(reg_weight_43_3), .partial_sum_in(reg_psum_43_3), .reg_activation(reg_activation_44_3), .reg_weight(reg_weight_44_3), .reg_partial_sum(reg_psum_44_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_4( .activation_in(reg_activation_44_3), .weight_in(reg_weight_43_4), .partial_sum_in(reg_psum_43_4), .reg_activation(reg_activation_44_4), .reg_weight(reg_weight_44_4), .reg_partial_sum(reg_psum_44_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_5( .activation_in(reg_activation_44_4), .weight_in(reg_weight_43_5), .partial_sum_in(reg_psum_43_5), .reg_activation(reg_activation_44_5), .reg_weight(reg_weight_44_5), .reg_partial_sum(reg_psum_44_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_6( .activation_in(reg_activation_44_5), .weight_in(reg_weight_43_6), .partial_sum_in(reg_psum_43_6), .reg_activation(reg_activation_44_6), .reg_weight(reg_weight_44_6), .reg_partial_sum(reg_psum_44_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_7( .activation_in(reg_activation_44_6), .weight_in(reg_weight_43_7), .partial_sum_in(reg_psum_43_7), .reg_activation(reg_activation_44_7), .reg_weight(reg_weight_44_7), .reg_partial_sum(reg_psum_44_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_8( .activation_in(reg_activation_44_7), .weight_in(reg_weight_43_8), .partial_sum_in(reg_psum_43_8), .reg_activation(reg_activation_44_8), .reg_weight(reg_weight_44_8), .reg_partial_sum(reg_psum_44_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_9( .activation_in(reg_activation_44_8), .weight_in(reg_weight_43_9), .partial_sum_in(reg_psum_43_9), .reg_activation(reg_activation_44_9), .reg_weight(reg_weight_44_9), .reg_partial_sum(reg_psum_44_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_10( .activation_in(reg_activation_44_9), .weight_in(reg_weight_43_10), .partial_sum_in(reg_psum_43_10), .reg_activation(reg_activation_44_10), .reg_weight(reg_weight_44_10), .reg_partial_sum(reg_psum_44_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_11( .activation_in(reg_activation_44_10), .weight_in(reg_weight_43_11), .partial_sum_in(reg_psum_43_11), .reg_activation(reg_activation_44_11), .reg_weight(reg_weight_44_11), .reg_partial_sum(reg_psum_44_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_12( .activation_in(reg_activation_44_11), .weight_in(reg_weight_43_12), .partial_sum_in(reg_psum_43_12), .reg_activation(reg_activation_44_12), .reg_weight(reg_weight_44_12), .reg_partial_sum(reg_psum_44_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_13( .activation_in(reg_activation_44_12), .weight_in(reg_weight_43_13), .partial_sum_in(reg_psum_43_13), .reg_activation(reg_activation_44_13), .reg_weight(reg_weight_44_13), .reg_partial_sum(reg_psum_44_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_14( .activation_in(reg_activation_44_13), .weight_in(reg_weight_43_14), .partial_sum_in(reg_psum_43_14), .reg_activation(reg_activation_44_14), .reg_weight(reg_weight_44_14), .reg_partial_sum(reg_psum_44_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_15( .activation_in(reg_activation_44_14), .weight_in(reg_weight_43_15), .partial_sum_in(reg_psum_43_15), .reg_activation(reg_activation_44_15), .reg_weight(reg_weight_44_15), .reg_partial_sum(reg_psum_44_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_16( .activation_in(reg_activation_44_15), .weight_in(reg_weight_43_16), .partial_sum_in(reg_psum_43_16), .reg_activation(reg_activation_44_16), .reg_weight(reg_weight_44_16), .reg_partial_sum(reg_psum_44_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_17( .activation_in(reg_activation_44_16), .weight_in(reg_weight_43_17), .partial_sum_in(reg_psum_43_17), .reg_activation(reg_activation_44_17), .reg_weight(reg_weight_44_17), .reg_partial_sum(reg_psum_44_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_18( .activation_in(reg_activation_44_17), .weight_in(reg_weight_43_18), .partial_sum_in(reg_psum_43_18), .reg_activation(reg_activation_44_18), .reg_weight(reg_weight_44_18), .reg_partial_sum(reg_psum_44_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_19( .activation_in(reg_activation_44_18), .weight_in(reg_weight_43_19), .partial_sum_in(reg_psum_43_19), .reg_activation(reg_activation_44_19), .reg_weight(reg_weight_44_19), .reg_partial_sum(reg_psum_44_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_20( .activation_in(reg_activation_44_19), .weight_in(reg_weight_43_20), .partial_sum_in(reg_psum_43_20), .reg_activation(reg_activation_44_20), .reg_weight(reg_weight_44_20), .reg_partial_sum(reg_psum_44_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_21( .activation_in(reg_activation_44_20), .weight_in(reg_weight_43_21), .partial_sum_in(reg_psum_43_21), .reg_activation(reg_activation_44_21), .reg_weight(reg_weight_44_21), .reg_partial_sum(reg_psum_44_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_22( .activation_in(reg_activation_44_21), .weight_in(reg_weight_43_22), .partial_sum_in(reg_psum_43_22), .reg_activation(reg_activation_44_22), .reg_weight(reg_weight_44_22), .reg_partial_sum(reg_psum_44_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_23( .activation_in(reg_activation_44_22), .weight_in(reg_weight_43_23), .partial_sum_in(reg_psum_43_23), .reg_activation(reg_activation_44_23), .reg_weight(reg_weight_44_23), .reg_partial_sum(reg_psum_44_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_24( .activation_in(reg_activation_44_23), .weight_in(reg_weight_43_24), .partial_sum_in(reg_psum_43_24), .reg_activation(reg_activation_44_24), .reg_weight(reg_weight_44_24), .reg_partial_sum(reg_psum_44_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_25( .activation_in(reg_activation_44_24), .weight_in(reg_weight_43_25), .partial_sum_in(reg_psum_43_25), .reg_activation(reg_activation_44_25), .reg_weight(reg_weight_44_25), .reg_partial_sum(reg_psum_44_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_26( .activation_in(reg_activation_44_25), .weight_in(reg_weight_43_26), .partial_sum_in(reg_psum_43_26), .reg_activation(reg_activation_44_26), .reg_weight(reg_weight_44_26), .reg_partial_sum(reg_psum_44_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_27( .activation_in(reg_activation_44_26), .weight_in(reg_weight_43_27), .partial_sum_in(reg_psum_43_27), .reg_activation(reg_activation_44_27), .reg_weight(reg_weight_44_27), .reg_partial_sum(reg_psum_44_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_28( .activation_in(reg_activation_44_27), .weight_in(reg_weight_43_28), .partial_sum_in(reg_psum_43_28), .reg_activation(reg_activation_44_28), .reg_weight(reg_weight_44_28), .reg_partial_sum(reg_psum_44_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_29( .activation_in(reg_activation_44_28), .weight_in(reg_weight_43_29), .partial_sum_in(reg_psum_43_29), .reg_activation(reg_activation_44_29), .reg_weight(reg_weight_44_29), .reg_partial_sum(reg_psum_44_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_30( .activation_in(reg_activation_44_29), .weight_in(reg_weight_43_30), .partial_sum_in(reg_psum_43_30), .reg_activation(reg_activation_44_30), .reg_weight(reg_weight_44_30), .reg_partial_sum(reg_psum_44_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_31( .activation_in(reg_activation_44_30), .weight_in(reg_weight_43_31), .partial_sum_in(reg_psum_43_31), .reg_activation(reg_activation_44_31), .reg_weight(reg_weight_44_31), .reg_partial_sum(reg_psum_44_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_32( .activation_in(reg_activation_44_31), .weight_in(reg_weight_43_32), .partial_sum_in(reg_psum_43_32), .reg_activation(reg_activation_44_32), .reg_weight(reg_weight_44_32), .reg_partial_sum(reg_psum_44_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_33( .activation_in(reg_activation_44_32), .weight_in(reg_weight_43_33), .partial_sum_in(reg_psum_43_33), .reg_activation(reg_activation_44_33), .reg_weight(reg_weight_44_33), .reg_partial_sum(reg_psum_44_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_34( .activation_in(reg_activation_44_33), .weight_in(reg_weight_43_34), .partial_sum_in(reg_psum_43_34), .reg_activation(reg_activation_44_34), .reg_weight(reg_weight_44_34), .reg_partial_sum(reg_psum_44_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_35( .activation_in(reg_activation_44_34), .weight_in(reg_weight_43_35), .partial_sum_in(reg_psum_43_35), .reg_activation(reg_activation_44_35), .reg_weight(reg_weight_44_35), .reg_partial_sum(reg_psum_44_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_36( .activation_in(reg_activation_44_35), .weight_in(reg_weight_43_36), .partial_sum_in(reg_psum_43_36), .reg_activation(reg_activation_44_36), .reg_weight(reg_weight_44_36), .reg_partial_sum(reg_psum_44_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_37( .activation_in(reg_activation_44_36), .weight_in(reg_weight_43_37), .partial_sum_in(reg_psum_43_37), .reg_activation(reg_activation_44_37), .reg_weight(reg_weight_44_37), .reg_partial_sum(reg_psum_44_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_38( .activation_in(reg_activation_44_37), .weight_in(reg_weight_43_38), .partial_sum_in(reg_psum_43_38), .reg_activation(reg_activation_44_38), .reg_weight(reg_weight_44_38), .reg_partial_sum(reg_psum_44_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_39( .activation_in(reg_activation_44_38), .weight_in(reg_weight_43_39), .partial_sum_in(reg_psum_43_39), .reg_activation(reg_activation_44_39), .reg_weight(reg_weight_44_39), .reg_partial_sum(reg_psum_44_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_40( .activation_in(reg_activation_44_39), .weight_in(reg_weight_43_40), .partial_sum_in(reg_psum_43_40), .reg_activation(reg_activation_44_40), .reg_weight(reg_weight_44_40), .reg_partial_sum(reg_psum_44_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_41( .activation_in(reg_activation_44_40), .weight_in(reg_weight_43_41), .partial_sum_in(reg_psum_43_41), .reg_activation(reg_activation_44_41), .reg_weight(reg_weight_44_41), .reg_partial_sum(reg_psum_44_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_42( .activation_in(reg_activation_44_41), .weight_in(reg_weight_43_42), .partial_sum_in(reg_psum_43_42), .reg_activation(reg_activation_44_42), .reg_weight(reg_weight_44_42), .reg_partial_sum(reg_psum_44_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_43( .activation_in(reg_activation_44_42), .weight_in(reg_weight_43_43), .partial_sum_in(reg_psum_43_43), .reg_activation(reg_activation_44_43), .reg_weight(reg_weight_44_43), .reg_partial_sum(reg_psum_44_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_44( .activation_in(reg_activation_44_43), .weight_in(reg_weight_43_44), .partial_sum_in(reg_psum_43_44), .reg_activation(reg_activation_44_44), .reg_weight(reg_weight_44_44), .reg_partial_sum(reg_psum_44_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_45( .activation_in(reg_activation_44_44), .weight_in(reg_weight_43_45), .partial_sum_in(reg_psum_43_45), .reg_activation(reg_activation_44_45), .reg_weight(reg_weight_44_45), .reg_partial_sum(reg_psum_44_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_46( .activation_in(reg_activation_44_45), .weight_in(reg_weight_43_46), .partial_sum_in(reg_psum_43_46), .reg_activation(reg_activation_44_46), .reg_weight(reg_weight_44_46), .reg_partial_sum(reg_psum_44_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_47( .activation_in(reg_activation_44_46), .weight_in(reg_weight_43_47), .partial_sum_in(reg_psum_43_47), .reg_activation(reg_activation_44_47), .reg_weight(reg_weight_44_47), .reg_partial_sum(reg_psum_44_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_48( .activation_in(reg_activation_44_47), .weight_in(reg_weight_43_48), .partial_sum_in(reg_psum_43_48), .reg_activation(reg_activation_44_48), .reg_weight(reg_weight_44_48), .reg_partial_sum(reg_psum_44_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_49( .activation_in(reg_activation_44_48), .weight_in(reg_weight_43_49), .partial_sum_in(reg_psum_43_49), .reg_activation(reg_activation_44_49), .reg_weight(reg_weight_44_49), .reg_partial_sum(reg_psum_44_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_50( .activation_in(reg_activation_44_49), .weight_in(reg_weight_43_50), .partial_sum_in(reg_psum_43_50), .reg_activation(reg_activation_44_50), .reg_weight(reg_weight_44_50), .reg_partial_sum(reg_psum_44_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_51( .activation_in(reg_activation_44_50), .weight_in(reg_weight_43_51), .partial_sum_in(reg_psum_43_51), .reg_activation(reg_activation_44_51), .reg_weight(reg_weight_44_51), .reg_partial_sum(reg_psum_44_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_52( .activation_in(reg_activation_44_51), .weight_in(reg_weight_43_52), .partial_sum_in(reg_psum_43_52), .reg_activation(reg_activation_44_52), .reg_weight(reg_weight_44_52), .reg_partial_sum(reg_psum_44_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_53( .activation_in(reg_activation_44_52), .weight_in(reg_weight_43_53), .partial_sum_in(reg_psum_43_53), .reg_activation(reg_activation_44_53), .reg_weight(reg_weight_44_53), .reg_partial_sum(reg_psum_44_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_54( .activation_in(reg_activation_44_53), .weight_in(reg_weight_43_54), .partial_sum_in(reg_psum_43_54), .reg_activation(reg_activation_44_54), .reg_weight(reg_weight_44_54), .reg_partial_sum(reg_psum_44_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_55( .activation_in(reg_activation_44_54), .weight_in(reg_weight_43_55), .partial_sum_in(reg_psum_43_55), .reg_activation(reg_activation_44_55), .reg_weight(reg_weight_44_55), .reg_partial_sum(reg_psum_44_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_56( .activation_in(reg_activation_44_55), .weight_in(reg_weight_43_56), .partial_sum_in(reg_psum_43_56), .reg_activation(reg_activation_44_56), .reg_weight(reg_weight_44_56), .reg_partial_sum(reg_psum_44_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_57( .activation_in(reg_activation_44_56), .weight_in(reg_weight_43_57), .partial_sum_in(reg_psum_43_57), .reg_activation(reg_activation_44_57), .reg_weight(reg_weight_44_57), .reg_partial_sum(reg_psum_44_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_58( .activation_in(reg_activation_44_57), .weight_in(reg_weight_43_58), .partial_sum_in(reg_psum_43_58), .reg_activation(reg_activation_44_58), .reg_weight(reg_weight_44_58), .reg_partial_sum(reg_psum_44_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_59( .activation_in(reg_activation_44_58), .weight_in(reg_weight_43_59), .partial_sum_in(reg_psum_43_59), .reg_activation(reg_activation_44_59), .reg_weight(reg_weight_44_59), .reg_partial_sum(reg_psum_44_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_60( .activation_in(reg_activation_44_59), .weight_in(reg_weight_43_60), .partial_sum_in(reg_psum_43_60), .reg_activation(reg_activation_44_60), .reg_weight(reg_weight_44_60), .reg_partial_sum(reg_psum_44_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_61( .activation_in(reg_activation_44_60), .weight_in(reg_weight_43_61), .partial_sum_in(reg_psum_43_61), .reg_activation(reg_activation_44_61), .reg_weight(reg_weight_44_61), .reg_partial_sum(reg_psum_44_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_62( .activation_in(reg_activation_44_61), .weight_in(reg_weight_43_62), .partial_sum_in(reg_psum_43_62), .reg_activation(reg_activation_44_62), .reg_weight(reg_weight_44_62), .reg_partial_sum(reg_psum_44_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U44_63( .activation_in(reg_activation_44_62), .weight_in(reg_weight_43_63), .partial_sum_in(reg_psum_43_63), .reg_weight(reg_weight_44_63), .reg_partial_sum(reg_psum_44_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_0( .activation_in(in_activation_45), .weight_in(reg_weight_44_0), .partial_sum_in(reg_psum_44_0), .reg_activation(reg_activation_45_0), .reg_weight(reg_weight_45_0), .reg_partial_sum(reg_psum_45_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_1( .activation_in(reg_activation_45_0), .weight_in(reg_weight_44_1), .partial_sum_in(reg_psum_44_1), .reg_activation(reg_activation_45_1), .reg_weight(reg_weight_45_1), .reg_partial_sum(reg_psum_45_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_2( .activation_in(reg_activation_45_1), .weight_in(reg_weight_44_2), .partial_sum_in(reg_psum_44_2), .reg_activation(reg_activation_45_2), .reg_weight(reg_weight_45_2), .reg_partial_sum(reg_psum_45_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_3( .activation_in(reg_activation_45_2), .weight_in(reg_weight_44_3), .partial_sum_in(reg_psum_44_3), .reg_activation(reg_activation_45_3), .reg_weight(reg_weight_45_3), .reg_partial_sum(reg_psum_45_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_4( .activation_in(reg_activation_45_3), .weight_in(reg_weight_44_4), .partial_sum_in(reg_psum_44_4), .reg_activation(reg_activation_45_4), .reg_weight(reg_weight_45_4), .reg_partial_sum(reg_psum_45_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_5( .activation_in(reg_activation_45_4), .weight_in(reg_weight_44_5), .partial_sum_in(reg_psum_44_5), .reg_activation(reg_activation_45_5), .reg_weight(reg_weight_45_5), .reg_partial_sum(reg_psum_45_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_6( .activation_in(reg_activation_45_5), .weight_in(reg_weight_44_6), .partial_sum_in(reg_psum_44_6), .reg_activation(reg_activation_45_6), .reg_weight(reg_weight_45_6), .reg_partial_sum(reg_psum_45_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_7( .activation_in(reg_activation_45_6), .weight_in(reg_weight_44_7), .partial_sum_in(reg_psum_44_7), .reg_activation(reg_activation_45_7), .reg_weight(reg_weight_45_7), .reg_partial_sum(reg_psum_45_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_8( .activation_in(reg_activation_45_7), .weight_in(reg_weight_44_8), .partial_sum_in(reg_psum_44_8), .reg_activation(reg_activation_45_8), .reg_weight(reg_weight_45_8), .reg_partial_sum(reg_psum_45_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_9( .activation_in(reg_activation_45_8), .weight_in(reg_weight_44_9), .partial_sum_in(reg_psum_44_9), .reg_activation(reg_activation_45_9), .reg_weight(reg_weight_45_9), .reg_partial_sum(reg_psum_45_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_10( .activation_in(reg_activation_45_9), .weight_in(reg_weight_44_10), .partial_sum_in(reg_psum_44_10), .reg_activation(reg_activation_45_10), .reg_weight(reg_weight_45_10), .reg_partial_sum(reg_psum_45_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_11( .activation_in(reg_activation_45_10), .weight_in(reg_weight_44_11), .partial_sum_in(reg_psum_44_11), .reg_activation(reg_activation_45_11), .reg_weight(reg_weight_45_11), .reg_partial_sum(reg_psum_45_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_12( .activation_in(reg_activation_45_11), .weight_in(reg_weight_44_12), .partial_sum_in(reg_psum_44_12), .reg_activation(reg_activation_45_12), .reg_weight(reg_weight_45_12), .reg_partial_sum(reg_psum_45_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_13( .activation_in(reg_activation_45_12), .weight_in(reg_weight_44_13), .partial_sum_in(reg_psum_44_13), .reg_activation(reg_activation_45_13), .reg_weight(reg_weight_45_13), .reg_partial_sum(reg_psum_45_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_14( .activation_in(reg_activation_45_13), .weight_in(reg_weight_44_14), .partial_sum_in(reg_psum_44_14), .reg_activation(reg_activation_45_14), .reg_weight(reg_weight_45_14), .reg_partial_sum(reg_psum_45_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_15( .activation_in(reg_activation_45_14), .weight_in(reg_weight_44_15), .partial_sum_in(reg_psum_44_15), .reg_activation(reg_activation_45_15), .reg_weight(reg_weight_45_15), .reg_partial_sum(reg_psum_45_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_16( .activation_in(reg_activation_45_15), .weight_in(reg_weight_44_16), .partial_sum_in(reg_psum_44_16), .reg_activation(reg_activation_45_16), .reg_weight(reg_weight_45_16), .reg_partial_sum(reg_psum_45_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_17( .activation_in(reg_activation_45_16), .weight_in(reg_weight_44_17), .partial_sum_in(reg_psum_44_17), .reg_activation(reg_activation_45_17), .reg_weight(reg_weight_45_17), .reg_partial_sum(reg_psum_45_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_18( .activation_in(reg_activation_45_17), .weight_in(reg_weight_44_18), .partial_sum_in(reg_psum_44_18), .reg_activation(reg_activation_45_18), .reg_weight(reg_weight_45_18), .reg_partial_sum(reg_psum_45_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_19( .activation_in(reg_activation_45_18), .weight_in(reg_weight_44_19), .partial_sum_in(reg_psum_44_19), .reg_activation(reg_activation_45_19), .reg_weight(reg_weight_45_19), .reg_partial_sum(reg_psum_45_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_20( .activation_in(reg_activation_45_19), .weight_in(reg_weight_44_20), .partial_sum_in(reg_psum_44_20), .reg_activation(reg_activation_45_20), .reg_weight(reg_weight_45_20), .reg_partial_sum(reg_psum_45_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_21( .activation_in(reg_activation_45_20), .weight_in(reg_weight_44_21), .partial_sum_in(reg_psum_44_21), .reg_activation(reg_activation_45_21), .reg_weight(reg_weight_45_21), .reg_partial_sum(reg_psum_45_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_22( .activation_in(reg_activation_45_21), .weight_in(reg_weight_44_22), .partial_sum_in(reg_psum_44_22), .reg_activation(reg_activation_45_22), .reg_weight(reg_weight_45_22), .reg_partial_sum(reg_psum_45_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_23( .activation_in(reg_activation_45_22), .weight_in(reg_weight_44_23), .partial_sum_in(reg_psum_44_23), .reg_activation(reg_activation_45_23), .reg_weight(reg_weight_45_23), .reg_partial_sum(reg_psum_45_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_24( .activation_in(reg_activation_45_23), .weight_in(reg_weight_44_24), .partial_sum_in(reg_psum_44_24), .reg_activation(reg_activation_45_24), .reg_weight(reg_weight_45_24), .reg_partial_sum(reg_psum_45_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_25( .activation_in(reg_activation_45_24), .weight_in(reg_weight_44_25), .partial_sum_in(reg_psum_44_25), .reg_activation(reg_activation_45_25), .reg_weight(reg_weight_45_25), .reg_partial_sum(reg_psum_45_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_26( .activation_in(reg_activation_45_25), .weight_in(reg_weight_44_26), .partial_sum_in(reg_psum_44_26), .reg_activation(reg_activation_45_26), .reg_weight(reg_weight_45_26), .reg_partial_sum(reg_psum_45_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_27( .activation_in(reg_activation_45_26), .weight_in(reg_weight_44_27), .partial_sum_in(reg_psum_44_27), .reg_activation(reg_activation_45_27), .reg_weight(reg_weight_45_27), .reg_partial_sum(reg_psum_45_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_28( .activation_in(reg_activation_45_27), .weight_in(reg_weight_44_28), .partial_sum_in(reg_psum_44_28), .reg_activation(reg_activation_45_28), .reg_weight(reg_weight_45_28), .reg_partial_sum(reg_psum_45_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_29( .activation_in(reg_activation_45_28), .weight_in(reg_weight_44_29), .partial_sum_in(reg_psum_44_29), .reg_activation(reg_activation_45_29), .reg_weight(reg_weight_45_29), .reg_partial_sum(reg_psum_45_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_30( .activation_in(reg_activation_45_29), .weight_in(reg_weight_44_30), .partial_sum_in(reg_psum_44_30), .reg_activation(reg_activation_45_30), .reg_weight(reg_weight_45_30), .reg_partial_sum(reg_psum_45_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_31( .activation_in(reg_activation_45_30), .weight_in(reg_weight_44_31), .partial_sum_in(reg_psum_44_31), .reg_activation(reg_activation_45_31), .reg_weight(reg_weight_45_31), .reg_partial_sum(reg_psum_45_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_32( .activation_in(reg_activation_45_31), .weight_in(reg_weight_44_32), .partial_sum_in(reg_psum_44_32), .reg_activation(reg_activation_45_32), .reg_weight(reg_weight_45_32), .reg_partial_sum(reg_psum_45_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_33( .activation_in(reg_activation_45_32), .weight_in(reg_weight_44_33), .partial_sum_in(reg_psum_44_33), .reg_activation(reg_activation_45_33), .reg_weight(reg_weight_45_33), .reg_partial_sum(reg_psum_45_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_34( .activation_in(reg_activation_45_33), .weight_in(reg_weight_44_34), .partial_sum_in(reg_psum_44_34), .reg_activation(reg_activation_45_34), .reg_weight(reg_weight_45_34), .reg_partial_sum(reg_psum_45_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_35( .activation_in(reg_activation_45_34), .weight_in(reg_weight_44_35), .partial_sum_in(reg_psum_44_35), .reg_activation(reg_activation_45_35), .reg_weight(reg_weight_45_35), .reg_partial_sum(reg_psum_45_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_36( .activation_in(reg_activation_45_35), .weight_in(reg_weight_44_36), .partial_sum_in(reg_psum_44_36), .reg_activation(reg_activation_45_36), .reg_weight(reg_weight_45_36), .reg_partial_sum(reg_psum_45_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_37( .activation_in(reg_activation_45_36), .weight_in(reg_weight_44_37), .partial_sum_in(reg_psum_44_37), .reg_activation(reg_activation_45_37), .reg_weight(reg_weight_45_37), .reg_partial_sum(reg_psum_45_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_38( .activation_in(reg_activation_45_37), .weight_in(reg_weight_44_38), .partial_sum_in(reg_psum_44_38), .reg_activation(reg_activation_45_38), .reg_weight(reg_weight_45_38), .reg_partial_sum(reg_psum_45_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_39( .activation_in(reg_activation_45_38), .weight_in(reg_weight_44_39), .partial_sum_in(reg_psum_44_39), .reg_activation(reg_activation_45_39), .reg_weight(reg_weight_45_39), .reg_partial_sum(reg_psum_45_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_40( .activation_in(reg_activation_45_39), .weight_in(reg_weight_44_40), .partial_sum_in(reg_psum_44_40), .reg_activation(reg_activation_45_40), .reg_weight(reg_weight_45_40), .reg_partial_sum(reg_psum_45_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_41( .activation_in(reg_activation_45_40), .weight_in(reg_weight_44_41), .partial_sum_in(reg_psum_44_41), .reg_activation(reg_activation_45_41), .reg_weight(reg_weight_45_41), .reg_partial_sum(reg_psum_45_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_42( .activation_in(reg_activation_45_41), .weight_in(reg_weight_44_42), .partial_sum_in(reg_psum_44_42), .reg_activation(reg_activation_45_42), .reg_weight(reg_weight_45_42), .reg_partial_sum(reg_psum_45_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_43( .activation_in(reg_activation_45_42), .weight_in(reg_weight_44_43), .partial_sum_in(reg_psum_44_43), .reg_activation(reg_activation_45_43), .reg_weight(reg_weight_45_43), .reg_partial_sum(reg_psum_45_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_44( .activation_in(reg_activation_45_43), .weight_in(reg_weight_44_44), .partial_sum_in(reg_psum_44_44), .reg_activation(reg_activation_45_44), .reg_weight(reg_weight_45_44), .reg_partial_sum(reg_psum_45_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_45( .activation_in(reg_activation_45_44), .weight_in(reg_weight_44_45), .partial_sum_in(reg_psum_44_45), .reg_activation(reg_activation_45_45), .reg_weight(reg_weight_45_45), .reg_partial_sum(reg_psum_45_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_46( .activation_in(reg_activation_45_45), .weight_in(reg_weight_44_46), .partial_sum_in(reg_psum_44_46), .reg_activation(reg_activation_45_46), .reg_weight(reg_weight_45_46), .reg_partial_sum(reg_psum_45_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_47( .activation_in(reg_activation_45_46), .weight_in(reg_weight_44_47), .partial_sum_in(reg_psum_44_47), .reg_activation(reg_activation_45_47), .reg_weight(reg_weight_45_47), .reg_partial_sum(reg_psum_45_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_48( .activation_in(reg_activation_45_47), .weight_in(reg_weight_44_48), .partial_sum_in(reg_psum_44_48), .reg_activation(reg_activation_45_48), .reg_weight(reg_weight_45_48), .reg_partial_sum(reg_psum_45_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_49( .activation_in(reg_activation_45_48), .weight_in(reg_weight_44_49), .partial_sum_in(reg_psum_44_49), .reg_activation(reg_activation_45_49), .reg_weight(reg_weight_45_49), .reg_partial_sum(reg_psum_45_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_50( .activation_in(reg_activation_45_49), .weight_in(reg_weight_44_50), .partial_sum_in(reg_psum_44_50), .reg_activation(reg_activation_45_50), .reg_weight(reg_weight_45_50), .reg_partial_sum(reg_psum_45_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_51( .activation_in(reg_activation_45_50), .weight_in(reg_weight_44_51), .partial_sum_in(reg_psum_44_51), .reg_activation(reg_activation_45_51), .reg_weight(reg_weight_45_51), .reg_partial_sum(reg_psum_45_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_52( .activation_in(reg_activation_45_51), .weight_in(reg_weight_44_52), .partial_sum_in(reg_psum_44_52), .reg_activation(reg_activation_45_52), .reg_weight(reg_weight_45_52), .reg_partial_sum(reg_psum_45_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_53( .activation_in(reg_activation_45_52), .weight_in(reg_weight_44_53), .partial_sum_in(reg_psum_44_53), .reg_activation(reg_activation_45_53), .reg_weight(reg_weight_45_53), .reg_partial_sum(reg_psum_45_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_54( .activation_in(reg_activation_45_53), .weight_in(reg_weight_44_54), .partial_sum_in(reg_psum_44_54), .reg_activation(reg_activation_45_54), .reg_weight(reg_weight_45_54), .reg_partial_sum(reg_psum_45_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_55( .activation_in(reg_activation_45_54), .weight_in(reg_weight_44_55), .partial_sum_in(reg_psum_44_55), .reg_activation(reg_activation_45_55), .reg_weight(reg_weight_45_55), .reg_partial_sum(reg_psum_45_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_56( .activation_in(reg_activation_45_55), .weight_in(reg_weight_44_56), .partial_sum_in(reg_psum_44_56), .reg_activation(reg_activation_45_56), .reg_weight(reg_weight_45_56), .reg_partial_sum(reg_psum_45_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_57( .activation_in(reg_activation_45_56), .weight_in(reg_weight_44_57), .partial_sum_in(reg_psum_44_57), .reg_activation(reg_activation_45_57), .reg_weight(reg_weight_45_57), .reg_partial_sum(reg_psum_45_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_58( .activation_in(reg_activation_45_57), .weight_in(reg_weight_44_58), .partial_sum_in(reg_psum_44_58), .reg_activation(reg_activation_45_58), .reg_weight(reg_weight_45_58), .reg_partial_sum(reg_psum_45_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_59( .activation_in(reg_activation_45_58), .weight_in(reg_weight_44_59), .partial_sum_in(reg_psum_44_59), .reg_activation(reg_activation_45_59), .reg_weight(reg_weight_45_59), .reg_partial_sum(reg_psum_45_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_60( .activation_in(reg_activation_45_59), .weight_in(reg_weight_44_60), .partial_sum_in(reg_psum_44_60), .reg_activation(reg_activation_45_60), .reg_weight(reg_weight_45_60), .reg_partial_sum(reg_psum_45_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_61( .activation_in(reg_activation_45_60), .weight_in(reg_weight_44_61), .partial_sum_in(reg_psum_44_61), .reg_activation(reg_activation_45_61), .reg_weight(reg_weight_45_61), .reg_partial_sum(reg_psum_45_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_62( .activation_in(reg_activation_45_61), .weight_in(reg_weight_44_62), .partial_sum_in(reg_psum_44_62), .reg_activation(reg_activation_45_62), .reg_weight(reg_weight_45_62), .reg_partial_sum(reg_psum_45_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U45_63( .activation_in(reg_activation_45_62), .weight_in(reg_weight_44_63), .partial_sum_in(reg_psum_44_63), .reg_weight(reg_weight_45_63), .reg_partial_sum(reg_psum_45_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_0( .activation_in(in_activation_46), .weight_in(reg_weight_45_0), .partial_sum_in(reg_psum_45_0), .reg_activation(reg_activation_46_0), .reg_weight(reg_weight_46_0), .reg_partial_sum(reg_psum_46_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_1( .activation_in(reg_activation_46_0), .weight_in(reg_weight_45_1), .partial_sum_in(reg_psum_45_1), .reg_activation(reg_activation_46_1), .reg_weight(reg_weight_46_1), .reg_partial_sum(reg_psum_46_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_2( .activation_in(reg_activation_46_1), .weight_in(reg_weight_45_2), .partial_sum_in(reg_psum_45_2), .reg_activation(reg_activation_46_2), .reg_weight(reg_weight_46_2), .reg_partial_sum(reg_psum_46_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_3( .activation_in(reg_activation_46_2), .weight_in(reg_weight_45_3), .partial_sum_in(reg_psum_45_3), .reg_activation(reg_activation_46_3), .reg_weight(reg_weight_46_3), .reg_partial_sum(reg_psum_46_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_4( .activation_in(reg_activation_46_3), .weight_in(reg_weight_45_4), .partial_sum_in(reg_psum_45_4), .reg_activation(reg_activation_46_4), .reg_weight(reg_weight_46_4), .reg_partial_sum(reg_psum_46_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_5( .activation_in(reg_activation_46_4), .weight_in(reg_weight_45_5), .partial_sum_in(reg_psum_45_5), .reg_activation(reg_activation_46_5), .reg_weight(reg_weight_46_5), .reg_partial_sum(reg_psum_46_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_6( .activation_in(reg_activation_46_5), .weight_in(reg_weight_45_6), .partial_sum_in(reg_psum_45_6), .reg_activation(reg_activation_46_6), .reg_weight(reg_weight_46_6), .reg_partial_sum(reg_psum_46_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_7( .activation_in(reg_activation_46_6), .weight_in(reg_weight_45_7), .partial_sum_in(reg_psum_45_7), .reg_activation(reg_activation_46_7), .reg_weight(reg_weight_46_7), .reg_partial_sum(reg_psum_46_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_8( .activation_in(reg_activation_46_7), .weight_in(reg_weight_45_8), .partial_sum_in(reg_psum_45_8), .reg_activation(reg_activation_46_8), .reg_weight(reg_weight_46_8), .reg_partial_sum(reg_psum_46_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_9( .activation_in(reg_activation_46_8), .weight_in(reg_weight_45_9), .partial_sum_in(reg_psum_45_9), .reg_activation(reg_activation_46_9), .reg_weight(reg_weight_46_9), .reg_partial_sum(reg_psum_46_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_10( .activation_in(reg_activation_46_9), .weight_in(reg_weight_45_10), .partial_sum_in(reg_psum_45_10), .reg_activation(reg_activation_46_10), .reg_weight(reg_weight_46_10), .reg_partial_sum(reg_psum_46_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_11( .activation_in(reg_activation_46_10), .weight_in(reg_weight_45_11), .partial_sum_in(reg_psum_45_11), .reg_activation(reg_activation_46_11), .reg_weight(reg_weight_46_11), .reg_partial_sum(reg_psum_46_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_12( .activation_in(reg_activation_46_11), .weight_in(reg_weight_45_12), .partial_sum_in(reg_psum_45_12), .reg_activation(reg_activation_46_12), .reg_weight(reg_weight_46_12), .reg_partial_sum(reg_psum_46_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_13( .activation_in(reg_activation_46_12), .weight_in(reg_weight_45_13), .partial_sum_in(reg_psum_45_13), .reg_activation(reg_activation_46_13), .reg_weight(reg_weight_46_13), .reg_partial_sum(reg_psum_46_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_14( .activation_in(reg_activation_46_13), .weight_in(reg_weight_45_14), .partial_sum_in(reg_psum_45_14), .reg_activation(reg_activation_46_14), .reg_weight(reg_weight_46_14), .reg_partial_sum(reg_psum_46_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_15( .activation_in(reg_activation_46_14), .weight_in(reg_weight_45_15), .partial_sum_in(reg_psum_45_15), .reg_activation(reg_activation_46_15), .reg_weight(reg_weight_46_15), .reg_partial_sum(reg_psum_46_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_16( .activation_in(reg_activation_46_15), .weight_in(reg_weight_45_16), .partial_sum_in(reg_psum_45_16), .reg_activation(reg_activation_46_16), .reg_weight(reg_weight_46_16), .reg_partial_sum(reg_psum_46_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_17( .activation_in(reg_activation_46_16), .weight_in(reg_weight_45_17), .partial_sum_in(reg_psum_45_17), .reg_activation(reg_activation_46_17), .reg_weight(reg_weight_46_17), .reg_partial_sum(reg_psum_46_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_18( .activation_in(reg_activation_46_17), .weight_in(reg_weight_45_18), .partial_sum_in(reg_psum_45_18), .reg_activation(reg_activation_46_18), .reg_weight(reg_weight_46_18), .reg_partial_sum(reg_psum_46_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_19( .activation_in(reg_activation_46_18), .weight_in(reg_weight_45_19), .partial_sum_in(reg_psum_45_19), .reg_activation(reg_activation_46_19), .reg_weight(reg_weight_46_19), .reg_partial_sum(reg_psum_46_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_20( .activation_in(reg_activation_46_19), .weight_in(reg_weight_45_20), .partial_sum_in(reg_psum_45_20), .reg_activation(reg_activation_46_20), .reg_weight(reg_weight_46_20), .reg_partial_sum(reg_psum_46_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_21( .activation_in(reg_activation_46_20), .weight_in(reg_weight_45_21), .partial_sum_in(reg_psum_45_21), .reg_activation(reg_activation_46_21), .reg_weight(reg_weight_46_21), .reg_partial_sum(reg_psum_46_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_22( .activation_in(reg_activation_46_21), .weight_in(reg_weight_45_22), .partial_sum_in(reg_psum_45_22), .reg_activation(reg_activation_46_22), .reg_weight(reg_weight_46_22), .reg_partial_sum(reg_psum_46_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_23( .activation_in(reg_activation_46_22), .weight_in(reg_weight_45_23), .partial_sum_in(reg_psum_45_23), .reg_activation(reg_activation_46_23), .reg_weight(reg_weight_46_23), .reg_partial_sum(reg_psum_46_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_24( .activation_in(reg_activation_46_23), .weight_in(reg_weight_45_24), .partial_sum_in(reg_psum_45_24), .reg_activation(reg_activation_46_24), .reg_weight(reg_weight_46_24), .reg_partial_sum(reg_psum_46_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_25( .activation_in(reg_activation_46_24), .weight_in(reg_weight_45_25), .partial_sum_in(reg_psum_45_25), .reg_activation(reg_activation_46_25), .reg_weight(reg_weight_46_25), .reg_partial_sum(reg_psum_46_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_26( .activation_in(reg_activation_46_25), .weight_in(reg_weight_45_26), .partial_sum_in(reg_psum_45_26), .reg_activation(reg_activation_46_26), .reg_weight(reg_weight_46_26), .reg_partial_sum(reg_psum_46_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_27( .activation_in(reg_activation_46_26), .weight_in(reg_weight_45_27), .partial_sum_in(reg_psum_45_27), .reg_activation(reg_activation_46_27), .reg_weight(reg_weight_46_27), .reg_partial_sum(reg_psum_46_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_28( .activation_in(reg_activation_46_27), .weight_in(reg_weight_45_28), .partial_sum_in(reg_psum_45_28), .reg_activation(reg_activation_46_28), .reg_weight(reg_weight_46_28), .reg_partial_sum(reg_psum_46_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_29( .activation_in(reg_activation_46_28), .weight_in(reg_weight_45_29), .partial_sum_in(reg_psum_45_29), .reg_activation(reg_activation_46_29), .reg_weight(reg_weight_46_29), .reg_partial_sum(reg_psum_46_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_30( .activation_in(reg_activation_46_29), .weight_in(reg_weight_45_30), .partial_sum_in(reg_psum_45_30), .reg_activation(reg_activation_46_30), .reg_weight(reg_weight_46_30), .reg_partial_sum(reg_psum_46_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_31( .activation_in(reg_activation_46_30), .weight_in(reg_weight_45_31), .partial_sum_in(reg_psum_45_31), .reg_activation(reg_activation_46_31), .reg_weight(reg_weight_46_31), .reg_partial_sum(reg_psum_46_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_32( .activation_in(reg_activation_46_31), .weight_in(reg_weight_45_32), .partial_sum_in(reg_psum_45_32), .reg_activation(reg_activation_46_32), .reg_weight(reg_weight_46_32), .reg_partial_sum(reg_psum_46_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_33( .activation_in(reg_activation_46_32), .weight_in(reg_weight_45_33), .partial_sum_in(reg_psum_45_33), .reg_activation(reg_activation_46_33), .reg_weight(reg_weight_46_33), .reg_partial_sum(reg_psum_46_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_34( .activation_in(reg_activation_46_33), .weight_in(reg_weight_45_34), .partial_sum_in(reg_psum_45_34), .reg_activation(reg_activation_46_34), .reg_weight(reg_weight_46_34), .reg_partial_sum(reg_psum_46_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_35( .activation_in(reg_activation_46_34), .weight_in(reg_weight_45_35), .partial_sum_in(reg_psum_45_35), .reg_activation(reg_activation_46_35), .reg_weight(reg_weight_46_35), .reg_partial_sum(reg_psum_46_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_36( .activation_in(reg_activation_46_35), .weight_in(reg_weight_45_36), .partial_sum_in(reg_psum_45_36), .reg_activation(reg_activation_46_36), .reg_weight(reg_weight_46_36), .reg_partial_sum(reg_psum_46_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_37( .activation_in(reg_activation_46_36), .weight_in(reg_weight_45_37), .partial_sum_in(reg_psum_45_37), .reg_activation(reg_activation_46_37), .reg_weight(reg_weight_46_37), .reg_partial_sum(reg_psum_46_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_38( .activation_in(reg_activation_46_37), .weight_in(reg_weight_45_38), .partial_sum_in(reg_psum_45_38), .reg_activation(reg_activation_46_38), .reg_weight(reg_weight_46_38), .reg_partial_sum(reg_psum_46_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_39( .activation_in(reg_activation_46_38), .weight_in(reg_weight_45_39), .partial_sum_in(reg_psum_45_39), .reg_activation(reg_activation_46_39), .reg_weight(reg_weight_46_39), .reg_partial_sum(reg_psum_46_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_40( .activation_in(reg_activation_46_39), .weight_in(reg_weight_45_40), .partial_sum_in(reg_psum_45_40), .reg_activation(reg_activation_46_40), .reg_weight(reg_weight_46_40), .reg_partial_sum(reg_psum_46_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_41( .activation_in(reg_activation_46_40), .weight_in(reg_weight_45_41), .partial_sum_in(reg_psum_45_41), .reg_activation(reg_activation_46_41), .reg_weight(reg_weight_46_41), .reg_partial_sum(reg_psum_46_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_42( .activation_in(reg_activation_46_41), .weight_in(reg_weight_45_42), .partial_sum_in(reg_psum_45_42), .reg_activation(reg_activation_46_42), .reg_weight(reg_weight_46_42), .reg_partial_sum(reg_psum_46_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_43( .activation_in(reg_activation_46_42), .weight_in(reg_weight_45_43), .partial_sum_in(reg_psum_45_43), .reg_activation(reg_activation_46_43), .reg_weight(reg_weight_46_43), .reg_partial_sum(reg_psum_46_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_44( .activation_in(reg_activation_46_43), .weight_in(reg_weight_45_44), .partial_sum_in(reg_psum_45_44), .reg_activation(reg_activation_46_44), .reg_weight(reg_weight_46_44), .reg_partial_sum(reg_psum_46_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_45( .activation_in(reg_activation_46_44), .weight_in(reg_weight_45_45), .partial_sum_in(reg_psum_45_45), .reg_activation(reg_activation_46_45), .reg_weight(reg_weight_46_45), .reg_partial_sum(reg_psum_46_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_46( .activation_in(reg_activation_46_45), .weight_in(reg_weight_45_46), .partial_sum_in(reg_psum_45_46), .reg_activation(reg_activation_46_46), .reg_weight(reg_weight_46_46), .reg_partial_sum(reg_psum_46_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_47( .activation_in(reg_activation_46_46), .weight_in(reg_weight_45_47), .partial_sum_in(reg_psum_45_47), .reg_activation(reg_activation_46_47), .reg_weight(reg_weight_46_47), .reg_partial_sum(reg_psum_46_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_48( .activation_in(reg_activation_46_47), .weight_in(reg_weight_45_48), .partial_sum_in(reg_psum_45_48), .reg_activation(reg_activation_46_48), .reg_weight(reg_weight_46_48), .reg_partial_sum(reg_psum_46_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_49( .activation_in(reg_activation_46_48), .weight_in(reg_weight_45_49), .partial_sum_in(reg_psum_45_49), .reg_activation(reg_activation_46_49), .reg_weight(reg_weight_46_49), .reg_partial_sum(reg_psum_46_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_50( .activation_in(reg_activation_46_49), .weight_in(reg_weight_45_50), .partial_sum_in(reg_psum_45_50), .reg_activation(reg_activation_46_50), .reg_weight(reg_weight_46_50), .reg_partial_sum(reg_psum_46_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_51( .activation_in(reg_activation_46_50), .weight_in(reg_weight_45_51), .partial_sum_in(reg_psum_45_51), .reg_activation(reg_activation_46_51), .reg_weight(reg_weight_46_51), .reg_partial_sum(reg_psum_46_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_52( .activation_in(reg_activation_46_51), .weight_in(reg_weight_45_52), .partial_sum_in(reg_psum_45_52), .reg_activation(reg_activation_46_52), .reg_weight(reg_weight_46_52), .reg_partial_sum(reg_psum_46_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_53( .activation_in(reg_activation_46_52), .weight_in(reg_weight_45_53), .partial_sum_in(reg_psum_45_53), .reg_activation(reg_activation_46_53), .reg_weight(reg_weight_46_53), .reg_partial_sum(reg_psum_46_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_54( .activation_in(reg_activation_46_53), .weight_in(reg_weight_45_54), .partial_sum_in(reg_psum_45_54), .reg_activation(reg_activation_46_54), .reg_weight(reg_weight_46_54), .reg_partial_sum(reg_psum_46_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_55( .activation_in(reg_activation_46_54), .weight_in(reg_weight_45_55), .partial_sum_in(reg_psum_45_55), .reg_activation(reg_activation_46_55), .reg_weight(reg_weight_46_55), .reg_partial_sum(reg_psum_46_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_56( .activation_in(reg_activation_46_55), .weight_in(reg_weight_45_56), .partial_sum_in(reg_psum_45_56), .reg_activation(reg_activation_46_56), .reg_weight(reg_weight_46_56), .reg_partial_sum(reg_psum_46_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_57( .activation_in(reg_activation_46_56), .weight_in(reg_weight_45_57), .partial_sum_in(reg_psum_45_57), .reg_activation(reg_activation_46_57), .reg_weight(reg_weight_46_57), .reg_partial_sum(reg_psum_46_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_58( .activation_in(reg_activation_46_57), .weight_in(reg_weight_45_58), .partial_sum_in(reg_psum_45_58), .reg_activation(reg_activation_46_58), .reg_weight(reg_weight_46_58), .reg_partial_sum(reg_psum_46_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_59( .activation_in(reg_activation_46_58), .weight_in(reg_weight_45_59), .partial_sum_in(reg_psum_45_59), .reg_activation(reg_activation_46_59), .reg_weight(reg_weight_46_59), .reg_partial_sum(reg_psum_46_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_60( .activation_in(reg_activation_46_59), .weight_in(reg_weight_45_60), .partial_sum_in(reg_psum_45_60), .reg_activation(reg_activation_46_60), .reg_weight(reg_weight_46_60), .reg_partial_sum(reg_psum_46_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_61( .activation_in(reg_activation_46_60), .weight_in(reg_weight_45_61), .partial_sum_in(reg_psum_45_61), .reg_activation(reg_activation_46_61), .reg_weight(reg_weight_46_61), .reg_partial_sum(reg_psum_46_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_62( .activation_in(reg_activation_46_61), .weight_in(reg_weight_45_62), .partial_sum_in(reg_psum_45_62), .reg_activation(reg_activation_46_62), .reg_weight(reg_weight_46_62), .reg_partial_sum(reg_psum_46_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U46_63( .activation_in(reg_activation_46_62), .weight_in(reg_weight_45_63), .partial_sum_in(reg_psum_45_63), .reg_weight(reg_weight_46_63), .reg_partial_sum(reg_psum_46_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_0( .activation_in(in_activation_47), .weight_in(reg_weight_46_0), .partial_sum_in(reg_psum_46_0), .reg_activation(reg_activation_47_0), .reg_weight(reg_weight_47_0), .reg_partial_sum(reg_psum_47_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_1( .activation_in(reg_activation_47_0), .weight_in(reg_weight_46_1), .partial_sum_in(reg_psum_46_1), .reg_activation(reg_activation_47_1), .reg_weight(reg_weight_47_1), .reg_partial_sum(reg_psum_47_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_2( .activation_in(reg_activation_47_1), .weight_in(reg_weight_46_2), .partial_sum_in(reg_psum_46_2), .reg_activation(reg_activation_47_2), .reg_weight(reg_weight_47_2), .reg_partial_sum(reg_psum_47_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_3( .activation_in(reg_activation_47_2), .weight_in(reg_weight_46_3), .partial_sum_in(reg_psum_46_3), .reg_activation(reg_activation_47_3), .reg_weight(reg_weight_47_3), .reg_partial_sum(reg_psum_47_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_4( .activation_in(reg_activation_47_3), .weight_in(reg_weight_46_4), .partial_sum_in(reg_psum_46_4), .reg_activation(reg_activation_47_4), .reg_weight(reg_weight_47_4), .reg_partial_sum(reg_psum_47_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_5( .activation_in(reg_activation_47_4), .weight_in(reg_weight_46_5), .partial_sum_in(reg_psum_46_5), .reg_activation(reg_activation_47_5), .reg_weight(reg_weight_47_5), .reg_partial_sum(reg_psum_47_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_6( .activation_in(reg_activation_47_5), .weight_in(reg_weight_46_6), .partial_sum_in(reg_psum_46_6), .reg_activation(reg_activation_47_6), .reg_weight(reg_weight_47_6), .reg_partial_sum(reg_psum_47_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_7( .activation_in(reg_activation_47_6), .weight_in(reg_weight_46_7), .partial_sum_in(reg_psum_46_7), .reg_activation(reg_activation_47_7), .reg_weight(reg_weight_47_7), .reg_partial_sum(reg_psum_47_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_8( .activation_in(reg_activation_47_7), .weight_in(reg_weight_46_8), .partial_sum_in(reg_psum_46_8), .reg_activation(reg_activation_47_8), .reg_weight(reg_weight_47_8), .reg_partial_sum(reg_psum_47_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_9( .activation_in(reg_activation_47_8), .weight_in(reg_weight_46_9), .partial_sum_in(reg_psum_46_9), .reg_activation(reg_activation_47_9), .reg_weight(reg_weight_47_9), .reg_partial_sum(reg_psum_47_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_10( .activation_in(reg_activation_47_9), .weight_in(reg_weight_46_10), .partial_sum_in(reg_psum_46_10), .reg_activation(reg_activation_47_10), .reg_weight(reg_weight_47_10), .reg_partial_sum(reg_psum_47_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_11( .activation_in(reg_activation_47_10), .weight_in(reg_weight_46_11), .partial_sum_in(reg_psum_46_11), .reg_activation(reg_activation_47_11), .reg_weight(reg_weight_47_11), .reg_partial_sum(reg_psum_47_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_12( .activation_in(reg_activation_47_11), .weight_in(reg_weight_46_12), .partial_sum_in(reg_psum_46_12), .reg_activation(reg_activation_47_12), .reg_weight(reg_weight_47_12), .reg_partial_sum(reg_psum_47_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_13( .activation_in(reg_activation_47_12), .weight_in(reg_weight_46_13), .partial_sum_in(reg_psum_46_13), .reg_activation(reg_activation_47_13), .reg_weight(reg_weight_47_13), .reg_partial_sum(reg_psum_47_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_14( .activation_in(reg_activation_47_13), .weight_in(reg_weight_46_14), .partial_sum_in(reg_psum_46_14), .reg_activation(reg_activation_47_14), .reg_weight(reg_weight_47_14), .reg_partial_sum(reg_psum_47_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_15( .activation_in(reg_activation_47_14), .weight_in(reg_weight_46_15), .partial_sum_in(reg_psum_46_15), .reg_activation(reg_activation_47_15), .reg_weight(reg_weight_47_15), .reg_partial_sum(reg_psum_47_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_16( .activation_in(reg_activation_47_15), .weight_in(reg_weight_46_16), .partial_sum_in(reg_psum_46_16), .reg_activation(reg_activation_47_16), .reg_weight(reg_weight_47_16), .reg_partial_sum(reg_psum_47_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_17( .activation_in(reg_activation_47_16), .weight_in(reg_weight_46_17), .partial_sum_in(reg_psum_46_17), .reg_activation(reg_activation_47_17), .reg_weight(reg_weight_47_17), .reg_partial_sum(reg_psum_47_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_18( .activation_in(reg_activation_47_17), .weight_in(reg_weight_46_18), .partial_sum_in(reg_psum_46_18), .reg_activation(reg_activation_47_18), .reg_weight(reg_weight_47_18), .reg_partial_sum(reg_psum_47_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_19( .activation_in(reg_activation_47_18), .weight_in(reg_weight_46_19), .partial_sum_in(reg_psum_46_19), .reg_activation(reg_activation_47_19), .reg_weight(reg_weight_47_19), .reg_partial_sum(reg_psum_47_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_20( .activation_in(reg_activation_47_19), .weight_in(reg_weight_46_20), .partial_sum_in(reg_psum_46_20), .reg_activation(reg_activation_47_20), .reg_weight(reg_weight_47_20), .reg_partial_sum(reg_psum_47_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_21( .activation_in(reg_activation_47_20), .weight_in(reg_weight_46_21), .partial_sum_in(reg_psum_46_21), .reg_activation(reg_activation_47_21), .reg_weight(reg_weight_47_21), .reg_partial_sum(reg_psum_47_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_22( .activation_in(reg_activation_47_21), .weight_in(reg_weight_46_22), .partial_sum_in(reg_psum_46_22), .reg_activation(reg_activation_47_22), .reg_weight(reg_weight_47_22), .reg_partial_sum(reg_psum_47_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_23( .activation_in(reg_activation_47_22), .weight_in(reg_weight_46_23), .partial_sum_in(reg_psum_46_23), .reg_activation(reg_activation_47_23), .reg_weight(reg_weight_47_23), .reg_partial_sum(reg_psum_47_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_24( .activation_in(reg_activation_47_23), .weight_in(reg_weight_46_24), .partial_sum_in(reg_psum_46_24), .reg_activation(reg_activation_47_24), .reg_weight(reg_weight_47_24), .reg_partial_sum(reg_psum_47_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_25( .activation_in(reg_activation_47_24), .weight_in(reg_weight_46_25), .partial_sum_in(reg_psum_46_25), .reg_activation(reg_activation_47_25), .reg_weight(reg_weight_47_25), .reg_partial_sum(reg_psum_47_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_26( .activation_in(reg_activation_47_25), .weight_in(reg_weight_46_26), .partial_sum_in(reg_psum_46_26), .reg_activation(reg_activation_47_26), .reg_weight(reg_weight_47_26), .reg_partial_sum(reg_psum_47_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_27( .activation_in(reg_activation_47_26), .weight_in(reg_weight_46_27), .partial_sum_in(reg_psum_46_27), .reg_activation(reg_activation_47_27), .reg_weight(reg_weight_47_27), .reg_partial_sum(reg_psum_47_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_28( .activation_in(reg_activation_47_27), .weight_in(reg_weight_46_28), .partial_sum_in(reg_psum_46_28), .reg_activation(reg_activation_47_28), .reg_weight(reg_weight_47_28), .reg_partial_sum(reg_psum_47_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_29( .activation_in(reg_activation_47_28), .weight_in(reg_weight_46_29), .partial_sum_in(reg_psum_46_29), .reg_activation(reg_activation_47_29), .reg_weight(reg_weight_47_29), .reg_partial_sum(reg_psum_47_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_30( .activation_in(reg_activation_47_29), .weight_in(reg_weight_46_30), .partial_sum_in(reg_psum_46_30), .reg_activation(reg_activation_47_30), .reg_weight(reg_weight_47_30), .reg_partial_sum(reg_psum_47_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_31( .activation_in(reg_activation_47_30), .weight_in(reg_weight_46_31), .partial_sum_in(reg_psum_46_31), .reg_activation(reg_activation_47_31), .reg_weight(reg_weight_47_31), .reg_partial_sum(reg_psum_47_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_32( .activation_in(reg_activation_47_31), .weight_in(reg_weight_46_32), .partial_sum_in(reg_psum_46_32), .reg_activation(reg_activation_47_32), .reg_weight(reg_weight_47_32), .reg_partial_sum(reg_psum_47_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_33( .activation_in(reg_activation_47_32), .weight_in(reg_weight_46_33), .partial_sum_in(reg_psum_46_33), .reg_activation(reg_activation_47_33), .reg_weight(reg_weight_47_33), .reg_partial_sum(reg_psum_47_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_34( .activation_in(reg_activation_47_33), .weight_in(reg_weight_46_34), .partial_sum_in(reg_psum_46_34), .reg_activation(reg_activation_47_34), .reg_weight(reg_weight_47_34), .reg_partial_sum(reg_psum_47_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_35( .activation_in(reg_activation_47_34), .weight_in(reg_weight_46_35), .partial_sum_in(reg_psum_46_35), .reg_activation(reg_activation_47_35), .reg_weight(reg_weight_47_35), .reg_partial_sum(reg_psum_47_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_36( .activation_in(reg_activation_47_35), .weight_in(reg_weight_46_36), .partial_sum_in(reg_psum_46_36), .reg_activation(reg_activation_47_36), .reg_weight(reg_weight_47_36), .reg_partial_sum(reg_psum_47_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_37( .activation_in(reg_activation_47_36), .weight_in(reg_weight_46_37), .partial_sum_in(reg_psum_46_37), .reg_activation(reg_activation_47_37), .reg_weight(reg_weight_47_37), .reg_partial_sum(reg_psum_47_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_38( .activation_in(reg_activation_47_37), .weight_in(reg_weight_46_38), .partial_sum_in(reg_psum_46_38), .reg_activation(reg_activation_47_38), .reg_weight(reg_weight_47_38), .reg_partial_sum(reg_psum_47_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_39( .activation_in(reg_activation_47_38), .weight_in(reg_weight_46_39), .partial_sum_in(reg_psum_46_39), .reg_activation(reg_activation_47_39), .reg_weight(reg_weight_47_39), .reg_partial_sum(reg_psum_47_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_40( .activation_in(reg_activation_47_39), .weight_in(reg_weight_46_40), .partial_sum_in(reg_psum_46_40), .reg_activation(reg_activation_47_40), .reg_weight(reg_weight_47_40), .reg_partial_sum(reg_psum_47_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_41( .activation_in(reg_activation_47_40), .weight_in(reg_weight_46_41), .partial_sum_in(reg_psum_46_41), .reg_activation(reg_activation_47_41), .reg_weight(reg_weight_47_41), .reg_partial_sum(reg_psum_47_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_42( .activation_in(reg_activation_47_41), .weight_in(reg_weight_46_42), .partial_sum_in(reg_psum_46_42), .reg_activation(reg_activation_47_42), .reg_weight(reg_weight_47_42), .reg_partial_sum(reg_psum_47_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_43( .activation_in(reg_activation_47_42), .weight_in(reg_weight_46_43), .partial_sum_in(reg_psum_46_43), .reg_activation(reg_activation_47_43), .reg_weight(reg_weight_47_43), .reg_partial_sum(reg_psum_47_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_44( .activation_in(reg_activation_47_43), .weight_in(reg_weight_46_44), .partial_sum_in(reg_psum_46_44), .reg_activation(reg_activation_47_44), .reg_weight(reg_weight_47_44), .reg_partial_sum(reg_psum_47_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_45( .activation_in(reg_activation_47_44), .weight_in(reg_weight_46_45), .partial_sum_in(reg_psum_46_45), .reg_activation(reg_activation_47_45), .reg_weight(reg_weight_47_45), .reg_partial_sum(reg_psum_47_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_46( .activation_in(reg_activation_47_45), .weight_in(reg_weight_46_46), .partial_sum_in(reg_psum_46_46), .reg_activation(reg_activation_47_46), .reg_weight(reg_weight_47_46), .reg_partial_sum(reg_psum_47_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_47( .activation_in(reg_activation_47_46), .weight_in(reg_weight_46_47), .partial_sum_in(reg_psum_46_47), .reg_activation(reg_activation_47_47), .reg_weight(reg_weight_47_47), .reg_partial_sum(reg_psum_47_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_48( .activation_in(reg_activation_47_47), .weight_in(reg_weight_46_48), .partial_sum_in(reg_psum_46_48), .reg_activation(reg_activation_47_48), .reg_weight(reg_weight_47_48), .reg_partial_sum(reg_psum_47_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_49( .activation_in(reg_activation_47_48), .weight_in(reg_weight_46_49), .partial_sum_in(reg_psum_46_49), .reg_activation(reg_activation_47_49), .reg_weight(reg_weight_47_49), .reg_partial_sum(reg_psum_47_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_50( .activation_in(reg_activation_47_49), .weight_in(reg_weight_46_50), .partial_sum_in(reg_psum_46_50), .reg_activation(reg_activation_47_50), .reg_weight(reg_weight_47_50), .reg_partial_sum(reg_psum_47_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_51( .activation_in(reg_activation_47_50), .weight_in(reg_weight_46_51), .partial_sum_in(reg_psum_46_51), .reg_activation(reg_activation_47_51), .reg_weight(reg_weight_47_51), .reg_partial_sum(reg_psum_47_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_52( .activation_in(reg_activation_47_51), .weight_in(reg_weight_46_52), .partial_sum_in(reg_psum_46_52), .reg_activation(reg_activation_47_52), .reg_weight(reg_weight_47_52), .reg_partial_sum(reg_psum_47_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_53( .activation_in(reg_activation_47_52), .weight_in(reg_weight_46_53), .partial_sum_in(reg_psum_46_53), .reg_activation(reg_activation_47_53), .reg_weight(reg_weight_47_53), .reg_partial_sum(reg_psum_47_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_54( .activation_in(reg_activation_47_53), .weight_in(reg_weight_46_54), .partial_sum_in(reg_psum_46_54), .reg_activation(reg_activation_47_54), .reg_weight(reg_weight_47_54), .reg_partial_sum(reg_psum_47_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_55( .activation_in(reg_activation_47_54), .weight_in(reg_weight_46_55), .partial_sum_in(reg_psum_46_55), .reg_activation(reg_activation_47_55), .reg_weight(reg_weight_47_55), .reg_partial_sum(reg_psum_47_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_56( .activation_in(reg_activation_47_55), .weight_in(reg_weight_46_56), .partial_sum_in(reg_psum_46_56), .reg_activation(reg_activation_47_56), .reg_weight(reg_weight_47_56), .reg_partial_sum(reg_psum_47_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_57( .activation_in(reg_activation_47_56), .weight_in(reg_weight_46_57), .partial_sum_in(reg_psum_46_57), .reg_activation(reg_activation_47_57), .reg_weight(reg_weight_47_57), .reg_partial_sum(reg_psum_47_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_58( .activation_in(reg_activation_47_57), .weight_in(reg_weight_46_58), .partial_sum_in(reg_psum_46_58), .reg_activation(reg_activation_47_58), .reg_weight(reg_weight_47_58), .reg_partial_sum(reg_psum_47_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_59( .activation_in(reg_activation_47_58), .weight_in(reg_weight_46_59), .partial_sum_in(reg_psum_46_59), .reg_activation(reg_activation_47_59), .reg_weight(reg_weight_47_59), .reg_partial_sum(reg_psum_47_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_60( .activation_in(reg_activation_47_59), .weight_in(reg_weight_46_60), .partial_sum_in(reg_psum_46_60), .reg_activation(reg_activation_47_60), .reg_weight(reg_weight_47_60), .reg_partial_sum(reg_psum_47_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_61( .activation_in(reg_activation_47_60), .weight_in(reg_weight_46_61), .partial_sum_in(reg_psum_46_61), .reg_activation(reg_activation_47_61), .reg_weight(reg_weight_47_61), .reg_partial_sum(reg_psum_47_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_62( .activation_in(reg_activation_47_61), .weight_in(reg_weight_46_62), .partial_sum_in(reg_psum_46_62), .reg_activation(reg_activation_47_62), .reg_weight(reg_weight_47_62), .reg_partial_sum(reg_psum_47_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U47_63( .activation_in(reg_activation_47_62), .weight_in(reg_weight_46_63), .partial_sum_in(reg_psum_46_63), .reg_weight(reg_weight_47_63), .reg_partial_sum(reg_psum_47_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_0( .activation_in(in_activation_48), .weight_in(reg_weight_47_0), .partial_sum_in(reg_psum_47_0), .reg_activation(reg_activation_48_0), .reg_weight(reg_weight_48_0), .reg_partial_sum(reg_psum_48_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_1( .activation_in(reg_activation_48_0), .weight_in(reg_weight_47_1), .partial_sum_in(reg_psum_47_1), .reg_activation(reg_activation_48_1), .reg_weight(reg_weight_48_1), .reg_partial_sum(reg_psum_48_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_2( .activation_in(reg_activation_48_1), .weight_in(reg_weight_47_2), .partial_sum_in(reg_psum_47_2), .reg_activation(reg_activation_48_2), .reg_weight(reg_weight_48_2), .reg_partial_sum(reg_psum_48_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_3( .activation_in(reg_activation_48_2), .weight_in(reg_weight_47_3), .partial_sum_in(reg_psum_47_3), .reg_activation(reg_activation_48_3), .reg_weight(reg_weight_48_3), .reg_partial_sum(reg_psum_48_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_4( .activation_in(reg_activation_48_3), .weight_in(reg_weight_47_4), .partial_sum_in(reg_psum_47_4), .reg_activation(reg_activation_48_4), .reg_weight(reg_weight_48_4), .reg_partial_sum(reg_psum_48_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_5( .activation_in(reg_activation_48_4), .weight_in(reg_weight_47_5), .partial_sum_in(reg_psum_47_5), .reg_activation(reg_activation_48_5), .reg_weight(reg_weight_48_5), .reg_partial_sum(reg_psum_48_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_6( .activation_in(reg_activation_48_5), .weight_in(reg_weight_47_6), .partial_sum_in(reg_psum_47_6), .reg_activation(reg_activation_48_6), .reg_weight(reg_weight_48_6), .reg_partial_sum(reg_psum_48_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_7( .activation_in(reg_activation_48_6), .weight_in(reg_weight_47_7), .partial_sum_in(reg_psum_47_7), .reg_activation(reg_activation_48_7), .reg_weight(reg_weight_48_7), .reg_partial_sum(reg_psum_48_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_8( .activation_in(reg_activation_48_7), .weight_in(reg_weight_47_8), .partial_sum_in(reg_psum_47_8), .reg_activation(reg_activation_48_8), .reg_weight(reg_weight_48_8), .reg_partial_sum(reg_psum_48_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_9( .activation_in(reg_activation_48_8), .weight_in(reg_weight_47_9), .partial_sum_in(reg_psum_47_9), .reg_activation(reg_activation_48_9), .reg_weight(reg_weight_48_9), .reg_partial_sum(reg_psum_48_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_10( .activation_in(reg_activation_48_9), .weight_in(reg_weight_47_10), .partial_sum_in(reg_psum_47_10), .reg_activation(reg_activation_48_10), .reg_weight(reg_weight_48_10), .reg_partial_sum(reg_psum_48_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_11( .activation_in(reg_activation_48_10), .weight_in(reg_weight_47_11), .partial_sum_in(reg_psum_47_11), .reg_activation(reg_activation_48_11), .reg_weight(reg_weight_48_11), .reg_partial_sum(reg_psum_48_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_12( .activation_in(reg_activation_48_11), .weight_in(reg_weight_47_12), .partial_sum_in(reg_psum_47_12), .reg_activation(reg_activation_48_12), .reg_weight(reg_weight_48_12), .reg_partial_sum(reg_psum_48_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_13( .activation_in(reg_activation_48_12), .weight_in(reg_weight_47_13), .partial_sum_in(reg_psum_47_13), .reg_activation(reg_activation_48_13), .reg_weight(reg_weight_48_13), .reg_partial_sum(reg_psum_48_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_14( .activation_in(reg_activation_48_13), .weight_in(reg_weight_47_14), .partial_sum_in(reg_psum_47_14), .reg_activation(reg_activation_48_14), .reg_weight(reg_weight_48_14), .reg_partial_sum(reg_psum_48_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_15( .activation_in(reg_activation_48_14), .weight_in(reg_weight_47_15), .partial_sum_in(reg_psum_47_15), .reg_activation(reg_activation_48_15), .reg_weight(reg_weight_48_15), .reg_partial_sum(reg_psum_48_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_16( .activation_in(reg_activation_48_15), .weight_in(reg_weight_47_16), .partial_sum_in(reg_psum_47_16), .reg_activation(reg_activation_48_16), .reg_weight(reg_weight_48_16), .reg_partial_sum(reg_psum_48_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_17( .activation_in(reg_activation_48_16), .weight_in(reg_weight_47_17), .partial_sum_in(reg_psum_47_17), .reg_activation(reg_activation_48_17), .reg_weight(reg_weight_48_17), .reg_partial_sum(reg_psum_48_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_18( .activation_in(reg_activation_48_17), .weight_in(reg_weight_47_18), .partial_sum_in(reg_psum_47_18), .reg_activation(reg_activation_48_18), .reg_weight(reg_weight_48_18), .reg_partial_sum(reg_psum_48_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_19( .activation_in(reg_activation_48_18), .weight_in(reg_weight_47_19), .partial_sum_in(reg_psum_47_19), .reg_activation(reg_activation_48_19), .reg_weight(reg_weight_48_19), .reg_partial_sum(reg_psum_48_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_20( .activation_in(reg_activation_48_19), .weight_in(reg_weight_47_20), .partial_sum_in(reg_psum_47_20), .reg_activation(reg_activation_48_20), .reg_weight(reg_weight_48_20), .reg_partial_sum(reg_psum_48_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_21( .activation_in(reg_activation_48_20), .weight_in(reg_weight_47_21), .partial_sum_in(reg_psum_47_21), .reg_activation(reg_activation_48_21), .reg_weight(reg_weight_48_21), .reg_partial_sum(reg_psum_48_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_22( .activation_in(reg_activation_48_21), .weight_in(reg_weight_47_22), .partial_sum_in(reg_psum_47_22), .reg_activation(reg_activation_48_22), .reg_weight(reg_weight_48_22), .reg_partial_sum(reg_psum_48_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_23( .activation_in(reg_activation_48_22), .weight_in(reg_weight_47_23), .partial_sum_in(reg_psum_47_23), .reg_activation(reg_activation_48_23), .reg_weight(reg_weight_48_23), .reg_partial_sum(reg_psum_48_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_24( .activation_in(reg_activation_48_23), .weight_in(reg_weight_47_24), .partial_sum_in(reg_psum_47_24), .reg_activation(reg_activation_48_24), .reg_weight(reg_weight_48_24), .reg_partial_sum(reg_psum_48_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_25( .activation_in(reg_activation_48_24), .weight_in(reg_weight_47_25), .partial_sum_in(reg_psum_47_25), .reg_activation(reg_activation_48_25), .reg_weight(reg_weight_48_25), .reg_partial_sum(reg_psum_48_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_26( .activation_in(reg_activation_48_25), .weight_in(reg_weight_47_26), .partial_sum_in(reg_psum_47_26), .reg_activation(reg_activation_48_26), .reg_weight(reg_weight_48_26), .reg_partial_sum(reg_psum_48_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_27( .activation_in(reg_activation_48_26), .weight_in(reg_weight_47_27), .partial_sum_in(reg_psum_47_27), .reg_activation(reg_activation_48_27), .reg_weight(reg_weight_48_27), .reg_partial_sum(reg_psum_48_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_28( .activation_in(reg_activation_48_27), .weight_in(reg_weight_47_28), .partial_sum_in(reg_psum_47_28), .reg_activation(reg_activation_48_28), .reg_weight(reg_weight_48_28), .reg_partial_sum(reg_psum_48_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_29( .activation_in(reg_activation_48_28), .weight_in(reg_weight_47_29), .partial_sum_in(reg_psum_47_29), .reg_activation(reg_activation_48_29), .reg_weight(reg_weight_48_29), .reg_partial_sum(reg_psum_48_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_30( .activation_in(reg_activation_48_29), .weight_in(reg_weight_47_30), .partial_sum_in(reg_psum_47_30), .reg_activation(reg_activation_48_30), .reg_weight(reg_weight_48_30), .reg_partial_sum(reg_psum_48_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_31( .activation_in(reg_activation_48_30), .weight_in(reg_weight_47_31), .partial_sum_in(reg_psum_47_31), .reg_activation(reg_activation_48_31), .reg_weight(reg_weight_48_31), .reg_partial_sum(reg_psum_48_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_32( .activation_in(reg_activation_48_31), .weight_in(reg_weight_47_32), .partial_sum_in(reg_psum_47_32), .reg_activation(reg_activation_48_32), .reg_weight(reg_weight_48_32), .reg_partial_sum(reg_psum_48_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_33( .activation_in(reg_activation_48_32), .weight_in(reg_weight_47_33), .partial_sum_in(reg_psum_47_33), .reg_activation(reg_activation_48_33), .reg_weight(reg_weight_48_33), .reg_partial_sum(reg_psum_48_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_34( .activation_in(reg_activation_48_33), .weight_in(reg_weight_47_34), .partial_sum_in(reg_psum_47_34), .reg_activation(reg_activation_48_34), .reg_weight(reg_weight_48_34), .reg_partial_sum(reg_psum_48_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_35( .activation_in(reg_activation_48_34), .weight_in(reg_weight_47_35), .partial_sum_in(reg_psum_47_35), .reg_activation(reg_activation_48_35), .reg_weight(reg_weight_48_35), .reg_partial_sum(reg_psum_48_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_36( .activation_in(reg_activation_48_35), .weight_in(reg_weight_47_36), .partial_sum_in(reg_psum_47_36), .reg_activation(reg_activation_48_36), .reg_weight(reg_weight_48_36), .reg_partial_sum(reg_psum_48_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_37( .activation_in(reg_activation_48_36), .weight_in(reg_weight_47_37), .partial_sum_in(reg_psum_47_37), .reg_activation(reg_activation_48_37), .reg_weight(reg_weight_48_37), .reg_partial_sum(reg_psum_48_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_38( .activation_in(reg_activation_48_37), .weight_in(reg_weight_47_38), .partial_sum_in(reg_psum_47_38), .reg_activation(reg_activation_48_38), .reg_weight(reg_weight_48_38), .reg_partial_sum(reg_psum_48_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_39( .activation_in(reg_activation_48_38), .weight_in(reg_weight_47_39), .partial_sum_in(reg_psum_47_39), .reg_activation(reg_activation_48_39), .reg_weight(reg_weight_48_39), .reg_partial_sum(reg_psum_48_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_40( .activation_in(reg_activation_48_39), .weight_in(reg_weight_47_40), .partial_sum_in(reg_psum_47_40), .reg_activation(reg_activation_48_40), .reg_weight(reg_weight_48_40), .reg_partial_sum(reg_psum_48_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_41( .activation_in(reg_activation_48_40), .weight_in(reg_weight_47_41), .partial_sum_in(reg_psum_47_41), .reg_activation(reg_activation_48_41), .reg_weight(reg_weight_48_41), .reg_partial_sum(reg_psum_48_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_42( .activation_in(reg_activation_48_41), .weight_in(reg_weight_47_42), .partial_sum_in(reg_psum_47_42), .reg_activation(reg_activation_48_42), .reg_weight(reg_weight_48_42), .reg_partial_sum(reg_psum_48_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_43( .activation_in(reg_activation_48_42), .weight_in(reg_weight_47_43), .partial_sum_in(reg_psum_47_43), .reg_activation(reg_activation_48_43), .reg_weight(reg_weight_48_43), .reg_partial_sum(reg_psum_48_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_44( .activation_in(reg_activation_48_43), .weight_in(reg_weight_47_44), .partial_sum_in(reg_psum_47_44), .reg_activation(reg_activation_48_44), .reg_weight(reg_weight_48_44), .reg_partial_sum(reg_psum_48_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_45( .activation_in(reg_activation_48_44), .weight_in(reg_weight_47_45), .partial_sum_in(reg_psum_47_45), .reg_activation(reg_activation_48_45), .reg_weight(reg_weight_48_45), .reg_partial_sum(reg_psum_48_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_46( .activation_in(reg_activation_48_45), .weight_in(reg_weight_47_46), .partial_sum_in(reg_psum_47_46), .reg_activation(reg_activation_48_46), .reg_weight(reg_weight_48_46), .reg_partial_sum(reg_psum_48_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_47( .activation_in(reg_activation_48_46), .weight_in(reg_weight_47_47), .partial_sum_in(reg_psum_47_47), .reg_activation(reg_activation_48_47), .reg_weight(reg_weight_48_47), .reg_partial_sum(reg_psum_48_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_48( .activation_in(reg_activation_48_47), .weight_in(reg_weight_47_48), .partial_sum_in(reg_psum_47_48), .reg_activation(reg_activation_48_48), .reg_weight(reg_weight_48_48), .reg_partial_sum(reg_psum_48_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_49( .activation_in(reg_activation_48_48), .weight_in(reg_weight_47_49), .partial_sum_in(reg_psum_47_49), .reg_activation(reg_activation_48_49), .reg_weight(reg_weight_48_49), .reg_partial_sum(reg_psum_48_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_50( .activation_in(reg_activation_48_49), .weight_in(reg_weight_47_50), .partial_sum_in(reg_psum_47_50), .reg_activation(reg_activation_48_50), .reg_weight(reg_weight_48_50), .reg_partial_sum(reg_psum_48_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_51( .activation_in(reg_activation_48_50), .weight_in(reg_weight_47_51), .partial_sum_in(reg_psum_47_51), .reg_activation(reg_activation_48_51), .reg_weight(reg_weight_48_51), .reg_partial_sum(reg_psum_48_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_52( .activation_in(reg_activation_48_51), .weight_in(reg_weight_47_52), .partial_sum_in(reg_psum_47_52), .reg_activation(reg_activation_48_52), .reg_weight(reg_weight_48_52), .reg_partial_sum(reg_psum_48_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_53( .activation_in(reg_activation_48_52), .weight_in(reg_weight_47_53), .partial_sum_in(reg_psum_47_53), .reg_activation(reg_activation_48_53), .reg_weight(reg_weight_48_53), .reg_partial_sum(reg_psum_48_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_54( .activation_in(reg_activation_48_53), .weight_in(reg_weight_47_54), .partial_sum_in(reg_psum_47_54), .reg_activation(reg_activation_48_54), .reg_weight(reg_weight_48_54), .reg_partial_sum(reg_psum_48_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_55( .activation_in(reg_activation_48_54), .weight_in(reg_weight_47_55), .partial_sum_in(reg_psum_47_55), .reg_activation(reg_activation_48_55), .reg_weight(reg_weight_48_55), .reg_partial_sum(reg_psum_48_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_56( .activation_in(reg_activation_48_55), .weight_in(reg_weight_47_56), .partial_sum_in(reg_psum_47_56), .reg_activation(reg_activation_48_56), .reg_weight(reg_weight_48_56), .reg_partial_sum(reg_psum_48_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_57( .activation_in(reg_activation_48_56), .weight_in(reg_weight_47_57), .partial_sum_in(reg_psum_47_57), .reg_activation(reg_activation_48_57), .reg_weight(reg_weight_48_57), .reg_partial_sum(reg_psum_48_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_58( .activation_in(reg_activation_48_57), .weight_in(reg_weight_47_58), .partial_sum_in(reg_psum_47_58), .reg_activation(reg_activation_48_58), .reg_weight(reg_weight_48_58), .reg_partial_sum(reg_psum_48_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_59( .activation_in(reg_activation_48_58), .weight_in(reg_weight_47_59), .partial_sum_in(reg_psum_47_59), .reg_activation(reg_activation_48_59), .reg_weight(reg_weight_48_59), .reg_partial_sum(reg_psum_48_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_60( .activation_in(reg_activation_48_59), .weight_in(reg_weight_47_60), .partial_sum_in(reg_psum_47_60), .reg_activation(reg_activation_48_60), .reg_weight(reg_weight_48_60), .reg_partial_sum(reg_psum_48_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_61( .activation_in(reg_activation_48_60), .weight_in(reg_weight_47_61), .partial_sum_in(reg_psum_47_61), .reg_activation(reg_activation_48_61), .reg_weight(reg_weight_48_61), .reg_partial_sum(reg_psum_48_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_62( .activation_in(reg_activation_48_61), .weight_in(reg_weight_47_62), .partial_sum_in(reg_psum_47_62), .reg_activation(reg_activation_48_62), .reg_weight(reg_weight_48_62), .reg_partial_sum(reg_psum_48_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U48_63( .activation_in(reg_activation_48_62), .weight_in(reg_weight_47_63), .partial_sum_in(reg_psum_47_63), .reg_weight(reg_weight_48_63), .reg_partial_sum(reg_psum_48_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_0( .activation_in(in_activation_49), .weight_in(reg_weight_48_0), .partial_sum_in(reg_psum_48_0), .reg_activation(reg_activation_49_0), .reg_weight(reg_weight_49_0), .reg_partial_sum(reg_psum_49_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_1( .activation_in(reg_activation_49_0), .weight_in(reg_weight_48_1), .partial_sum_in(reg_psum_48_1), .reg_activation(reg_activation_49_1), .reg_weight(reg_weight_49_1), .reg_partial_sum(reg_psum_49_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_2( .activation_in(reg_activation_49_1), .weight_in(reg_weight_48_2), .partial_sum_in(reg_psum_48_2), .reg_activation(reg_activation_49_2), .reg_weight(reg_weight_49_2), .reg_partial_sum(reg_psum_49_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_3( .activation_in(reg_activation_49_2), .weight_in(reg_weight_48_3), .partial_sum_in(reg_psum_48_3), .reg_activation(reg_activation_49_3), .reg_weight(reg_weight_49_3), .reg_partial_sum(reg_psum_49_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_4( .activation_in(reg_activation_49_3), .weight_in(reg_weight_48_4), .partial_sum_in(reg_psum_48_4), .reg_activation(reg_activation_49_4), .reg_weight(reg_weight_49_4), .reg_partial_sum(reg_psum_49_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_5( .activation_in(reg_activation_49_4), .weight_in(reg_weight_48_5), .partial_sum_in(reg_psum_48_5), .reg_activation(reg_activation_49_5), .reg_weight(reg_weight_49_5), .reg_partial_sum(reg_psum_49_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_6( .activation_in(reg_activation_49_5), .weight_in(reg_weight_48_6), .partial_sum_in(reg_psum_48_6), .reg_activation(reg_activation_49_6), .reg_weight(reg_weight_49_6), .reg_partial_sum(reg_psum_49_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_7( .activation_in(reg_activation_49_6), .weight_in(reg_weight_48_7), .partial_sum_in(reg_psum_48_7), .reg_activation(reg_activation_49_7), .reg_weight(reg_weight_49_7), .reg_partial_sum(reg_psum_49_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_8( .activation_in(reg_activation_49_7), .weight_in(reg_weight_48_8), .partial_sum_in(reg_psum_48_8), .reg_activation(reg_activation_49_8), .reg_weight(reg_weight_49_8), .reg_partial_sum(reg_psum_49_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_9( .activation_in(reg_activation_49_8), .weight_in(reg_weight_48_9), .partial_sum_in(reg_psum_48_9), .reg_activation(reg_activation_49_9), .reg_weight(reg_weight_49_9), .reg_partial_sum(reg_psum_49_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_10( .activation_in(reg_activation_49_9), .weight_in(reg_weight_48_10), .partial_sum_in(reg_psum_48_10), .reg_activation(reg_activation_49_10), .reg_weight(reg_weight_49_10), .reg_partial_sum(reg_psum_49_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_11( .activation_in(reg_activation_49_10), .weight_in(reg_weight_48_11), .partial_sum_in(reg_psum_48_11), .reg_activation(reg_activation_49_11), .reg_weight(reg_weight_49_11), .reg_partial_sum(reg_psum_49_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_12( .activation_in(reg_activation_49_11), .weight_in(reg_weight_48_12), .partial_sum_in(reg_psum_48_12), .reg_activation(reg_activation_49_12), .reg_weight(reg_weight_49_12), .reg_partial_sum(reg_psum_49_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_13( .activation_in(reg_activation_49_12), .weight_in(reg_weight_48_13), .partial_sum_in(reg_psum_48_13), .reg_activation(reg_activation_49_13), .reg_weight(reg_weight_49_13), .reg_partial_sum(reg_psum_49_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_14( .activation_in(reg_activation_49_13), .weight_in(reg_weight_48_14), .partial_sum_in(reg_psum_48_14), .reg_activation(reg_activation_49_14), .reg_weight(reg_weight_49_14), .reg_partial_sum(reg_psum_49_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_15( .activation_in(reg_activation_49_14), .weight_in(reg_weight_48_15), .partial_sum_in(reg_psum_48_15), .reg_activation(reg_activation_49_15), .reg_weight(reg_weight_49_15), .reg_partial_sum(reg_psum_49_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_16( .activation_in(reg_activation_49_15), .weight_in(reg_weight_48_16), .partial_sum_in(reg_psum_48_16), .reg_activation(reg_activation_49_16), .reg_weight(reg_weight_49_16), .reg_partial_sum(reg_psum_49_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_17( .activation_in(reg_activation_49_16), .weight_in(reg_weight_48_17), .partial_sum_in(reg_psum_48_17), .reg_activation(reg_activation_49_17), .reg_weight(reg_weight_49_17), .reg_partial_sum(reg_psum_49_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_18( .activation_in(reg_activation_49_17), .weight_in(reg_weight_48_18), .partial_sum_in(reg_psum_48_18), .reg_activation(reg_activation_49_18), .reg_weight(reg_weight_49_18), .reg_partial_sum(reg_psum_49_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_19( .activation_in(reg_activation_49_18), .weight_in(reg_weight_48_19), .partial_sum_in(reg_psum_48_19), .reg_activation(reg_activation_49_19), .reg_weight(reg_weight_49_19), .reg_partial_sum(reg_psum_49_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_20( .activation_in(reg_activation_49_19), .weight_in(reg_weight_48_20), .partial_sum_in(reg_psum_48_20), .reg_activation(reg_activation_49_20), .reg_weight(reg_weight_49_20), .reg_partial_sum(reg_psum_49_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_21( .activation_in(reg_activation_49_20), .weight_in(reg_weight_48_21), .partial_sum_in(reg_psum_48_21), .reg_activation(reg_activation_49_21), .reg_weight(reg_weight_49_21), .reg_partial_sum(reg_psum_49_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_22( .activation_in(reg_activation_49_21), .weight_in(reg_weight_48_22), .partial_sum_in(reg_psum_48_22), .reg_activation(reg_activation_49_22), .reg_weight(reg_weight_49_22), .reg_partial_sum(reg_psum_49_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_23( .activation_in(reg_activation_49_22), .weight_in(reg_weight_48_23), .partial_sum_in(reg_psum_48_23), .reg_activation(reg_activation_49_23), .reg_weight(reg_weight_49_23), .reg_partial_sum(reg_psum_49_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_24( .activation_in(reg_activation_49_23), .weight_in(reg_weight_48_24), .partial_sum_in(reg_psum_48_24), .reg_activation(reg_activation_49_24), .reg_weight(reg_weight_49_24), .reg_partial_sum(reg_psum_49_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_25( .activation_in(reg_activation_49_24), .weight_in(reg_weight_48_25), .partial_sum_in(reg_psum_48_25), .reg_activation(reg_activation_49_25), .reg_weight(reg_weight_49_25), .reg_partial_sum(reg_psum_49_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_26( .activation_in(reg_activation_49_25), .weight_in(reg_weight_48_26), .partial_sum_in(reg_psum_48_26), .reg_activation(reg_activation_49_26), .reg_weight(reg_weight_49_26), .reg_partial_sum(reg_psum_49_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_27( .activation_in(reg_activation_49_26), .weight_in(reg_weight_48_27), .partial_sum_in(reg_psum_48_27), .reg_activation(reg_activation_49_27), .reg_weight(reg_weight_49_27), .reg_partial_sum(reg_psum_49_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_28( .activation_in(reg_activation_49_27), .weight_in(reg_weight_48_28), .partial_sum_in(reg_psum_48_28), .reg_activation(reg_activation_49_28), .reg_weight(reg_weight_49_28), .reg_partial_sum(reg_psum_49_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_29( .activation_in(reg_activation_49_28), .weight_in(reg_weight_48_29), .partial_sum_in(reg_psum_48_29), .reg_activation(reg_activation_49_29), .reg_weight(reg_weight_49_29), .reg_partial_sum(reg_psum_49_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_30( .activation_in(reg_activation_49_29), .weight_in(reg_weight_48_30), .partial_sum_in(reg_psum_48_30), .reg_activation(reg_activation_49_30), .reg_weight(reg_weight_49_30), .reg_partial_sum(reg_psum_49_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_31( .activation_in(reg_activation_49_30), .weight_in(reg_weight_48_31), .partial_sum_in(reg_psum_48_31), .reg_activation(reg_activation_49_31), .reg_weight(reg_weight_49_31), .reg_partial_sum(reg_psum_49_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_32( .activation_in(reg_activation_49_31), .weight_in(reg_weight_48_32), .partial_sum_in(reg_psum_48_32), .reg_activation(reg_activation_49_32), .reg_weight(reg_weight_49_32), .reg_partial_sum(reg_psum_49_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_33( .activation_in(reg_activation_49_32), .weight_in(reg_weight_48_33), .partial_sum_in(reg_psum_48_33), .reg_activation(reg_activation_49_33), .reg_weight(reg_weight_49_33), .reg_partial_sum(reg_psum_49_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_34( .activation_in(reg_activation_49_33), .weight_in(reg_weight_48_34), .partial_sum_in(reg_psum_48_34), .reg_activation(reg_activation_49_34), .reg_weight(reg_weight_49_34), .reg_partial_sum(reg_psum_49_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_35( .activation_in(reg_activation_49_34), .weight_in(reg_weight_48_35), .partial_sum_in(reg_psum_48_35), .reg_activation(reg_activation_49_35), .reg_weight(reg_weight_49_35), .reg_partial_sum(reg_psum_49_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_36( .activation_in(reg_activation_49_35), .weight_in(reg_weight_48_36), .partial_sum_in(reg_psum_48_36), .reg_activation(reg_activation_49_36), .reg_weight(reg_weight_49_36), .reg_partial_sum(reg_psum_49_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_37( .activation_in(reg_activation_49_36), .weight_in(reg_weight_48_37), .partial_sum_in(reg_psum_48_37), .reg_activation(reg_activation_49_37), .reg_weight(reg_weight_49_37), .reg_partial_sum(reg_psum_49_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_38( .activation_in(reg_activation_49_37), .weight_in(reg_weight_48_38), .partial_sum_in(reg_psum_48_38), .reg_activation(reg_activation_49_38), .reg_weight(reg_weight_49_38), .reg_partial_sum(reg_psum_49_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_39( .activation_in(reg_activation_49_38), .weight_in(reg_weight_48_39), .partial_sum_in(reg_psum_48_39), .reg_activation(reg_activation_49_39), .reg_weight(reg_weight_49_39), .reg_partial_sum(reg_psum_49_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_40( .activation_in(reg_activation_49_39), .weight_in(reg_weight_48_40), .partial_sum_in(reg_psum_48_40), .reg_activation(reg_activation_49_40), .reg_weight(reg_weight_49_40), .reg_partial_sum(reg_psum_49_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_41( .activation_in(reg_activation_49_40), .weight_in(reg_weight_48_41), .partial_sum_in(reg_psum_48_41), .reg_activation(reg_activation_49_41), .reg_weight(reg_weight_49_41), .reg_partial_sum(reg_psum_49_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_42( .activation_in(reg_activation_49_41), .weight_in(reg_weight_48_42), .partial_sum_in(reg_psum_48_42), .reg_activation(reg_activation_49_42), .reg_weight(reg_weight_49_42), .reg_partial_sum(reg_psum_49_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_43( .activation_in(reg_activation_49_42), .weight_in(reg_weight_48_43), .partial_sum_in(reg_psum_48_43), .reg_activation(reg_activation_49_43), .reg_weight(reg_weight_49_43), .reg_partial_sum(reg_psum_49_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_44( .activation_in(reg_activation_49_43), .weight_in(reg_weight_48_44), .partial_sum_in(reg_psum_48_44), .reg_activation(reg_activation_49_44), .reg_weight(reg_weight_49_44), .reg_partial_sum(reg_psum_49_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_45( .activation_in(reg_activation_49_44), .weight_in(reg_weight_48_45), .partial_sum_in(reg_psum_48_45), .reg_activation(reg_activation_49_45), .reg_weight(reg_weight_49_45), .reg_partial_sum(reg_psum_49_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_46( .activation_in(reg_activation_49_45), .weight_in(reg_weight_48_46), .partial_sum_in(reg_psum_48_46), .reg_activation(reg_activation_49_46), .reg_weight(reg_weight_49_46), .reg_partial_sum(reg_psum_49_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_47( .activation_in(reg_activation_49_46), .weight_in(reg_weight_48_47), .partial_sum_in(reg_psum_48_47), .reg_activation(reg_activation_49_47), .reg_weight(reg_weight_49_47), .reg_partial_sum(reg_psum_49_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_48( .activation_in(reg_activation_49_47), .weight_in(reg_weight_48_48), .partial_sum_in(reg_psum_48_48), .reg_activation(reg_activation_49_48), .reg_weight(reg_weight_49_48), .reg_partial_sum(reg_psum_49_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_49( .activation_in(reg_activation_49_48), .weight_in(reg_weight_48_49), .partial_sum_in(reg_psum_48_49), .reg_activation(reg_activation_49_49), .reg_weight(reg_weight_49_49), .reg_partial_sum(reg_psum_49_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_50( .activation_in(reg_activation_49_49), .weight_in(reg_weight_48_50), .partial_sum_in(reg_psum_48_50), .reg_activation(reg_activation_49_50), .reg_weight(reg_weight_49_50), .reg_partial_sum(reg_psum_49_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_51( .activation_in(reg_activation_49_50), .weight_in(reg_weight_48_51), .partial_sum_in(reg_psum_48_51), .reg_activation(reg_activation_49_51), .reg_weight(reg_weight_49_51), .reg_partial_sum(reg_psum_49_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_52( .activation_in(reg_activation_49_51), .weight_in(reg_weight_48_52), .partial_sum_in(reg_psum_48_52), .reg_activation(reg_activation_49_52), .reg_weight(reg_weight_49_52), .reg_partial_sum(reg_psum_49_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_53( .activation_in(reg_activation_49_52), .weight_in(reg_weight_48_53), .partial_sum_in(reg_psum_48_53), .reg_activation(reg_activation_49_53), .reg_weight(reg_weight_49_53), .reg_partial_sum(reg_psum_49_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_54( .activation_in(reg_activation_49_53), .weight_in(reg_weight_48_54), .partial_sum_in(reg_psum_48_54), .reg_activation(reg_activation_49_54), .reg_weight(reg_weight_49_54), .reg_partial_sum(reg_psum_49_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_55( .activation_in(reg_activation_49_54), .weight_in(reg_weight_48_55), .partial_sum_in(reg_psum_48_55), .reg_activation(reg_activation_49_55), .reg_weight(reg_weight_49_55), .reg_partial_sum(reg_psum_49_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_56( .activation_in(reg_activation_49_55), .weight_in(reg_weight_48_56), .partial_sum_in(reg_psum_48_56), .reg_activation(reg_activation_49_56), .reg_weight(reg_weight_49_56), .reg_partial_sum(reg_psum_49_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_57( .activation_in(reg_activation_49_56), .weight_in(reg_weight_48_57), .partial_sum_in(reg_psum_48_57), .reg_activation(reg_activation_49_57), .reg_weight(reg_weight_49_57), .reg_partial_sum(reg_psum_49_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_58( .activation_in(reg_activation_49_57), .weight_in(reg_weight_48_58), .partial_sum_in(reg_psum_48_58), .reg_activation(reg_activation_49_58), .reg_weight(reg_weight_49_58), .reg_partial_sum(reg_psum_49_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_59( .activation_in(reg_activation_49_58), .weight_in(reg_weight_48_59), .partial_sum_in(reg_psum_48_59), .reg_activation(reg_activation_49_59), .reg_weight(reg_weight_49_59), .reg_partial_sum(reg_psum_49_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_60( .activation_in(reg_activation_49_59), .weight_in(reg_weight_48_60), .partial_sum_in(reg_psum_48_60), .reg_activation(reg_activation_49_60), .reg_weight(reg_weight_49_60), .reg_partial_sum(reg_psum_49_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_61( .activation_in(reg_activation_49_60), .weight_in(reg_weight_48_61), .partial_sum_in(reg_psum_48_61), .reg_activation(reg_activation_49_61), .reg_weight(reg_weight_49_61), .reg_partial_sum(reg_psum_49_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_62( .activation_in(reg_activation_49_61), .weight_in(reg_weight_48_62), .partial_sum_in(reg_psum_48_62), .reg_activation(reg_activation_49_62), .reg_weight(reg_weight_49_62), .reg_partial_sum(reg_psum_49_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U49_63( .activation_in(reg_activation_49_62), .weight_in(reg_weight_48_63), .partial_sum_in(reg_psum_48_63), .reg_weight(reg_weight_49_63), .reg_partial_sum(reg_psum_49_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_0( .activation_in(in_activation_50), .weight_in(reg_weight_49_0), .partial_sum_in(reg_psum_49_0), .reg_activation(reg_activation_50_0), .reg_weight(reg_weight_50_0), .reg_partial_sum(reg_psum_50_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_1( .activation_in(reg_activation_50_0), .weight_in(reg_weight_49_1), .partial_sum_in(reg_psum_49_1), .reg_activation(reg_activation_50_1), .reg_weight(reg_weight_50_1), .reg_partial_sum(reg_psum_50_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_2( .activation_in(reg_activation_50_1), .weight_in(reg_weight_49_2), .partial_sum_in(reg_psum_49_2), .reg_activation(reg_activation_50_2), .reg_weight(reg_weight_50_2), .reg_partial_sum(reg_psum_50_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_3( .activation_in(reg_activation_50_2), .weight_in(reg_weight_49_3), .partial_sum_in(reg_psum_49_3), .reg_activation(reg_activation_50_3), .reg_weight(reg_weight_50_3), .reg_partial_sum(reg_psum_50_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_4( .activation_in(reg_activation_50_3), .weight_in(reg_weight_49_4), .partial_sum_in(reg_psum_49_4), .reg_activation(reg_activation_50_4), .reg_weight(reg_weight_50_4), .reg_partial_sum(reg_psum_50_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_5( .activation_in(reg_activation_50_4), .weight_in(reg_weight_49_5), .partial_sum_in(reg_psum_49_5), .reg_activation(reg_activation_50_5), .reg_weight(reg_weight_50_5), .reg_partial_sum(reg_psum_50_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_6( .activation_in(reg_activation_50_5), .weight_in(reg_weight_49_6), .partial_sum_in(reg_psum_49_6), .reg_activation(reg_activation_50_6), .reg_weight(reg_weight_50_6), .reg_partial_sum(reg_psum_50_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_7( .activation_in(reg_activation_50_6), .weight_in(reg_weight_49_7), .partial_sum_in(reg_psum_49_7), .reg_activation(reg_activation_50_7), .reg_weight(reg_weight_50_7), .reg_partial_sum(reg_psum_50_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_8( .activation_in(reg_activation_50_7), .weight_in(reg_weight_49_8), .partial_sum_in(reg_psum_49_8), .reg_activation(reg_activation_50_8), .reg_weight(reg_weight_50_8), .reg_partial_sum(reg_psum_50_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_9( .activation_in(reg_activation_50_8), .weight_in(reg_weight_49_9), .partial_sum_in(reg_psum_49_9), .reg_activation(reg_activation_50_9), .reg_weight(reg_weight_50_9), .reg_partial_sum(reg_psum_50_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_10( .activation_in(reg_activation_50_9), .weight_in(reg_weight_49_10), .partial_sum_in(reg_psum_49_10), .reg_activation(reg_activation_50_10), .reg_weight(reg_weight_50_10), .reg_partial_sum(reg_psum_50_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_11( .activation_in(reg_activation_50_10), .weight_in(reg_weight_49_11), .partial_sum_in(reg_psum_49_11), .reg_activation(reg_activation_50_11), .reg_weight(reg_weight_50_11), .reg_partial_sum(reg_psum_50_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_12( .activation_in(reg_activation_50_11), .weight_in(reg_weight_49_12), .partial_sum_in(reg_psum_49_12), .reg_activation(reg_activation_50_12), .reg_weight(reg_weight_50_12), .reg_partial_sum(reg_psum_50_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_13( .activation_in(reg_activation_50_12), .weight_in(reg_weight_49_13), .partial_sum_in(reg_psum_49_13), .reg_activation(reg_activation_50_13), .reg_weight(reg_weight_50_13), .reg_partial_sum(reg_psum_50_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_14( .activation_in(reg_activation_50_13), .weight_in(reg_weight_49_14), .partial_sum_in(reg_psum_49_14), .reg_activation(reg_activation_50_14), .reg_weight(reg_weight_50_14), .reg_partial_sum(reg_psum_50_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_15( .activation_in(reg_activation_50_14), .weight_in(reg_weight_49_15), .partial_sum_in(reg_psum_49_15), .reg_activation(reg_activation_50_15), .reg_weight(reg_weight_50_15), .reg_partial_sum(reg_psum_50_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_16( .activation_in(reg_activation_50_15), .weight_in(reg_weight_49_16), .partial_sum_in(reg_psum_49_16), .reg_activation(reg_activation_50_16), .reg_weight(reg_weight_50_16), .reg_partial_sum(reg_psum_50_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_17( .activation_in(reg_activation_50_16), .weight_in(reg_weight_49_17), .partial_sum_in(reg_psum_49_17), .reg_activation(reg_activation_50_17), .reg_weight(reg_weight_50_17), .reg_partial_sum(reg_psum_50_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_18( .activation_in(reg_activation_50_17), .weight_in(reg_weight_49_18), .partial_sum_in(reg_psum_49_18), .reg_activation(reg_activation_50_18), .reg_weight(reg_weight_50_18), .reg_partial_sum(reg_psum_50_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_19( .activation_in(reg_activation_50_18), .weight_in(reg_weight_49_19), .partial_sum_in(reg_psum_49_19), .reg_activation(reg_activation_50_19), .reg_weight(reg_weight_50_19), .reg_partial_sum(reg_psum_50_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_20( .activation_in(reg_activation_50_19), .weight_in(reg_weight_49_20), .partial_sum_in(reg_psum_49_20), .reg_activation(reg_activation_50_20), .reg_weight(reg_weight_50_20), .reg_partial_sum(reg_psum_50_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_21( .activation_in(reg_activation_50_20), .weight_in(reg_weight_49_21), .partial_sum_in(reg_psum_49_21), .reg_activation(reg_activation_50_21), .reg_weight(reg_weight_50_21), .reg_partial_sum(reg_psum_50_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_22( .activation_in(reg_activation_50_21), .weight_in(reg_weight_49_22), .partial_sum_in(reg_psum_49_22), .reg_activation(reg_activation_50_22), .reg_weight(reg_weight_50_22), .reg_partial_sum(reg_psum_50_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_23( .activation_in(reg_activation_50_22), .weight_in(reg_weight_49_23), .partial_sum_in(reg_psum_49_23), .reg_activation(reg_activation_50_23), .reg_weight(reg_weight_50_23), .reg_partial_sum(reg_psum_50_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_24( .activation_in(reg_activation_50_23), .weight_in(reg_weight_49_24), .partial_sum_in(reg_psum_49_24), .reg_activation(reg_activation_50_24), .reg_weight(reg_weight_50_24), .reg_partial_sum(reg_psum_50_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_25( .activation_in(reg_activation_50_24), .weight_in(reg_weight_49_25), .partial_sum_in(reg_psum_49_25), .reg_activation(reg_activation_50_25), .reg_weight(reg_weight_50_25), .reg_partial_sum(reg_psum_50_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_26( .activation_in(reg_activation_50_25), .weight_in(reg_weight_49_26), .partial_sum_in(reg_psum_49_26), .reg_activation(reg_activation_50_26), .reg_weight(reg_weight_50_26), .reg_partial_sum(reg_psum_50_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_27( .activation_in(reg_activation_50_26), .weight_in(reg_weight_49_27), .partial_sum_in(reg_psum_49_27), .reg_activation(reg_activation_50_27), .reg_weight(reg_weight_50_27), .reg_partial_sum(reg_psum_50_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_28( .activation_in(reg_activation_50_27), .weight_in(reg_weight_49_28), .partial_sum_in(reg_psum_49_28), .reg_activation(reg_activation_50_28), .reg_weight(reg_weight_50_28), .reg_partial_sum(reg_psum_50_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_29( .activation_in(reg_activation_50_28), .weight_in(reg_weight_49_29), .partial_sum_in(reg_psum_49_29), .reg_activation(reg_activation_50_29), .reg_weight(reg_weight_50_29), .reg_partial_sum(reg_psum_50_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_30( .activation_in(reg_activation_50_29), .weight_in(reg_weight_49_30), .partial_sum_in(reg_psum_49_30), .reg_activation(reg_activation_50_30), .reg_weight(reg_weight_50_30), .reg_partial_sum(reg_psum_50_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_31( .activation_in(reg_activation_50_30), .weight_in(reg_weight_49_31), .partial_sum_in(reg_psum_49_31), .reg_activation(reg_activation_50_31), .reg_weight(reg_weight_50_31), .reg_partial_sum(reg_psum_50_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_32( .activation_in(reg_activation_50_31), .weight_in(reg_weight_49_32), .partial_sum_in(reg_psum_49_32), .reg_activation(reg_activation_50_32), .reg_weight(reg_weight_50_32), .reg_partial_sum(reg_psum_50_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_33( .activation_in(reg_activation_50_32), .weight_in(reg_weight_49_33), .partial_sum_in(reg_psum_49_33), .reg_activation(reg_activation_50_33), .reg_weight(reg_weight_50_33), .reg_partial_sum(reg_psum_50_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_34( .activation_in(reg_activation_50_33), .weight_in(reg_weight_49_34), .partial_sum_in(reg_psum_49_34), .reg_activation(reg_activation_50_34), .reg_weight(reg_weight_50_34), .reg_partial_sum(reg_psum_50_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_35( .activation_in(reg_activation_50_34), .weight_in(reg_weight_49_35), .partial_sum_in(reg_psum_49_35), .reg_activation(reg_activation_50_35), .reg_weight(reg_weight_50_35), .reg_partial_sum(reg_psum_50_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_36( .activation_in(reg_activation_50_35), .weight_in(reg_weight_49_36), .partial_sum_in(reg_psum_49_36), .reg_activation(reg_activation_50_36), .reg_weight(reg_weight_50_36), .reg_partial_sum(reg_psum_50_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_37( .activation_in(reg_activation_50_36), .weight_in(reg_weight_49_37), .partial_sum_in(reg_psum_49_37), .reg_activation(reg_activation_50_37), .reg_weight(reg_weight_50_37), .reg_partial_sum(reg_psum_50_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_38( .activation_in(reg_activation_50_37), .weight_in(reg_weight_49_38), .partial_sum_in(reg_psum_49_38), .reg_activation(reg_activation_50_38), .reg_weight(reg_weight_50_38), .reg_partial_sum(reg_psum_50_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_39( .activation_in(reg_activation_50_38), .weight_in(reg_weight_49_39), .partial_sum_in(reg_psum_49_39), .reg_activation(reg_activation_50_39), .reg_weight(reg_weight_50_39), .reg_partial_sum(reg_psum_50_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_40( .activation_in(reg_activation_50_39), .weight_in(reg_weight_49_40), .partial_sum_in(reg_psum_49_40), .reg_activation(reg_activation_50_40), .reg_weight(reg_weight_50_40), .reg_partial_sum(reg_psum_50_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_41( .activation_in(reg_activation_50_40), .weight_in(reg_weight_49_41), .partial_sum_in(reg_psum_49_41), .reg_activation(reg_activation_50_41), .reg_weight(reg_weight_50_41), .reg_partial_sum(reg_psum_50_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_42( .activation_in(reg_activation_50_41), .weight_in(reg_weight_49_42), .partial_sum_in(reg_psum_49_42), .reg_activation(reg_activation_50_42), .reg_weight(reg_weight_50_42), .reg_partial_sum(reg_psum_50_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_43( .activation_in(reg_activation_50_42), .weight_in(reg_weight_49_43), .partial_sum_in(reg_psum_49_43), .reg_activation(reg_activation_50_43), .reg_weight(reg_weight_50_43), .reg_partial_sum(reg_psum_50_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_44( .activation_in(reg_activation_50_43), .weight_in(reg_weight_49_44), .partial_sum_in(reg_psum_49_44), .reg_activation(reg_activation_50_44), .reg_weight(reg_weight_50_44), .reg_partial_sum(reg_psum_50_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_45( .activation_in(reg_activation_50_44), .weight_in(reg_weight_49_45), .partial_sum_in(reg_psum_49_45), .reg_activation(reg_activation_50_45), .reg_weight(reg_weight_50_45), .reg_partial_sum(reg_psum_50_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_46( .activation_in(reg_activation_50_45), .weight_in(reg_weight_49_46), .partial_sum_in(reg_psum_49_46), .reg_activation(reg_activation_50_46), .reg_weight(reg_weight_50_46), .reg_partial_sum(reg_psum_50_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_47( .activation_in(reg_activation_50_46), .weight_in(reg_weight_49_47), .partial_sum_in(reg_psum_49_47), .reg_activation(reg_activation_50_47), .reg_weight(reg_weight_50_47), .reg_partial_sum(reg_psum_50_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_48( .activation_in(reg_activation_50_47), .weight_in(reg_weight_49_48), .partial_sum_in(reg_psum_49_48), .reg_activation(reg_activation_50_48), .reg_weight(reg_weight_50_48), .reg_partial_sum(reg_psum_50_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_49( .activation_in(reg_activation_50_48), .weight_in(reg_weight_49_49), .partial_sum_in(reg_psum_49_49), .reg_activation(reg_activation_50_49), .reg_weight(reg_weight_50_49), .reg_partial_sum(reg_psum_50_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_50( .activation_in(reg_activation_50_49), .weight_in(reg_weight_49_50), .partial_sum_in(reg_psum_49_50), .reg_activation(reg_activation_50_50), .reg_weight(reg_weight_50_50), .reg_partial_sum(reg_psum_50_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_51( .activation_in(reg_activation_50_50), .weight_in(reg_weight_49_51), .partial_sum_in(reg_psum_49_51), .reg_activation(reg_activation_50_51), .reg_weight(reg_weight_50_51), .reg_partial_sum(reg_psum_50_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_52( .activation_in(reg_activation_50_51), .weight_in(reg_weight_49_52), .partial_sum_in(reg_psum_49_52), .reg_activation(reg_activation_50_52), .reg_weight(reg_weight_50_52), .reg_partial_sum(reg_psum_50_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_53( .activation_in(reg_activation_50_52), .weight_in(reg_weight_49_53), .partial_sum_in(reg_psum_49_53), .reg_activation(reg_activation_50_53), .reg_weight(reg_weight_50_53), .reg_partial_sum(reg_psum_50_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_54( .activation_in(reg_activation_50_53), .weight_in(reg_weight_49_54), .partial_sum_in(reg_psum_49_54), .reg_activation(reg_activation_50_54), .reg_weight(reg_weight_50_54), .reg_partial_sum(reg_psum_50_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_55( .activation_in(reg_activation_50_54), .weight_in(reg_weight_49_55), .partial_sum_in(reg_psum_49_55), .reg_activation(reg_activation_50_55), .reg_weight(reg_weight_50_55), .reg_partial_sum(reg_psum_50_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_56( .activation_in(reg_activation_50_55), .weight_in(reg_weight_49_56), .partial_sum_in(reg_psum_49_56), .reg_activation(reg_activation_50_56), .reg_weight(reg_weight_50_56), .reg_partial_sum(reg_psum_50_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_57( .activation_in(reg_activation_50_56), .weight_in(reg_weight_49_57), .partial_sum_in(reg_psum_49_57), .reg_activation(reg_activation_50_57), .reg_weight(reg_weight_50_57), .reg_partial_sum(reg_psum_50_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_58( .activation_in(reg_activation_50_57), .weight_in(reg_weight_49_58), .partial_sum_in(reg_psum_49_58), .reg_activation(reg_activation_50_58), .reg_weight(reg_weight_50_58), .reg_partial_sum(reg_psum_50_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_59( .activation_in(reg_activation_50_58), .weight_in(reg_weight_49_59), .partial_sum_in(reg_psum_49_59), .reg_activation(reg_activation_50_59), .reg_weight(reg_weight_50_59), .reg_partial_sum(reg_psum_50_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_60( .activation_in(reg_activation_50_59), .weight_in(reg_weight_49_60), .partial_sum_in(reg_psum_49_60), .reg_activation(reg_activation_50_60), .reg_weight(reg_weight_50_60), .reg_partial_sum(reg_psum_50_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_61( .activation_in(reg_activation_50_60), .weight_in(reg_weight_49_61), .partial_sum_in(reg_psum_49_61), .reg_activation(reg_activation_50_61), .reg_weight(reg_weight_50_61), .reg_partial_sum(reg_psum_50_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_62( .activation_in(reg_activation_50_61), .weight_in(reg_weight_49_62), .partial_sum_in(reg_psum_49_62), .reg_activation(reg_activation_50_62), .reg_weight(reg_weight_50_62), .reg_partial_sum(reg_psum_50_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U50_63( .activation_in(reg_activation_50_62), .weight_in(reg_weight_49_63), .partial_sum_in(reg_psum_49_63), .reg_weight(reg_weight_50_63), .reg_partial_sum(reg_psum_50_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_0( .activation_in(in_activation_51), .weight_in(reg_weight_50_0), .partial_sum_in(reg_psum_50_0), .reg_activation(reg_activation_51_0), .reg_weight(reg_weight_51_0), .reg_partial_sum(reg_psum_51_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_1( .activation_in(reg_activation_51_0), .weight_in(reg_weight_50_1), .partial_sum_in(reg_psum_50_1), .reg_activation(reg_activation_51_1), .reg_weight(reg_weight_51_1), .reg_partial_sum(reg_psum_51_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_2( .activation_in(reg_activation_51_1), .weight_in(reg_weight_50_2), .partial_sum_in(reg_psum_50_2), .reg_activation(reg_activation_51_2), .reg_weight(reg_weight_51_2), .reg_partial_sum(reg_psum_51_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_3( .activation_in(reg_activation_51_2), .weight_in(reg_weight_50_3), .partial_sum_in(reg_psum_50_3), .reg_activation(reg_activation_51_3), .reg_weight(reg_weight_51_3), .reg_partial_sum(reg_psum_51_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_4( .activation_in(reg_activation_51_3), .weight_in(reg_weight_50_4), .partial_sum_in(reg_psum_50_4), .reg_activation(reg_activation_51_4), .reg_weight(reg_weight_51_4), .reg_partial_sum(reg_psum_51_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_5( .activation_in(reg_activation_51_4), .weight_in(reg_weight_50_5), .partial_sum_in(reg_psum_50_5), .reg_activation(reg_activation_51_5), .reg_weight(reg_weight_51_5), .reg_partial_sum(reg_psum_51_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_6( .activation_in(reg_activation_51_5), .weight_in(reg_weight_50_6), .partial_sum_in(reg_psum_50_6), .reg_activation(reg_activation_51_6), .reg_weight(reg_weight_51_6), .reg_partial_sum(reg_psum_51_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_7( .activation_in(reg_activation_51_6), .weight_in(reg_weight_50_7), .partial_sum_in(reg_psum_50_7), .reg_activation(reg_activation_51_7), .reg_weight(reg_weight_51_7), .reg_partial_sum(reg_psum_51_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_8( .activation_in(reg_activation_51_7), .weight_in(reg_weight_50_8), .partial_sum_in(reg_psum_50_8), .reg_activation(reg_activation_51_8), .reg_weight(reg_weight_51_8), .reg_partial_sum(reg_psum_51_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_9( .activation_in(reg_activation_51_8), .weight_in(reg_weight_50_9), .partial_sum_in(reg_psum_50_9), .reg_activation(reg_activation_51_9), .reg_weight(reg_weight_51_9), .reg_partial_sum(reg_psum_51_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_10( .activation_in(reg_activation_51_9), .weight_in(reg_weight_50_10), .partial_sum_in(reg_psum_50_10), .reg_activation(reg_activation_51_10), .reg_weight(reg_weight_51_10), .reg_partial_sum(reg_psum_51_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_11( .activation_in(reg_activation_51_10), .weight_in(reg_weight_50_11), .partial_sum_in(reg_psum_50_11), .reg_activation(reg_activation_51_11), .reg_weight(reg_weight_51_11), .reg_partial_sum(reg_psum_51_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_12( .activation_in(reg_activation_51_11), .weight_in(reg_weight_50_12), .partial_sum_in(reg_psum_50_12), .reg_activation(reg_activation_51_12), .reg_weight(reg_weight_51_12), .reg_partial_sum(reg_psum_51_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_13( .activation_in(reg_activation_51_12), .weight_in(reg_weight_50_13), .partial_sum_in(reg_psum_50_13), .reg_activation(reg_activation_51_13), .reg_weight(reg_weight_51_13), .reg_partial_sum(reg_psum_51_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_14( .activation_in(reg_activation_51_13), .weight_in(reg_weight_50_14), .partial_sum_in(reg_psum_50_14), .reg_activation(reg_activation_51_14), .reg_weight(reg_weight_51_14), .reg_partial_sum(reg_psum_51_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_15( .activation_in(reg_activation_51_14), .weight_in(reg_weight_50_15), .partial_sum_in(reg_psum_50_15), .reg_activation(reg_activation_51_15), .reg_weight(reg_weight_51_15), .reg_partial_sum(reg_psum_51_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_16( .activation_in(reg_activation_51_15), .weight_in(reg_weight_50_16), .partial_sum_in(reg_psum_50_16), .reg_activation(reg_activation_51_16), .reg_weight(reg_weight_51_16), .reg_partial_sum(reg_psum_51_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_17( .activation_in(reg_activation_51_16), .weight_in(reg_weight_50_17), .partial_sum_in(reg_psum_50_17), .reg_activation(reg_activation_51_17), .reg_weight(reg_weight_51_17), .reg_partial_sum(reg_psum_51_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_18( .activation_in(reg_activation_51_17), .weight_in(reg_weight_50_18), .partial_sum_in(reg_psum_50_18), .reg_activation(reg_activation_51_18), .reg_weight(reg_weight_51_18), .reg_partial_sum(reg_psum_51_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_19( .activation_in(reg_activation_51_18), .weight_in(reg_weight_50_19), .partial_sum_in(reg_psum_50_19), .reg_activation(reg_activation_51_19), .reg_weight(reg_weight_51_19), .reg_partial_sum(reg_psum_51_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_20( .activation_in(reg_activation_51_19), .weight_in(reg_weight_50_20), .partial_sum_in(reg_psum_50_20), .reg_activation(reg_activation_51_20), .reg_weight(reg_weight_51_20), .reg_partial_sum(reg_psum_51_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_21( .activation_in(reg_activation_51_20), .weight_in(reg_weight_50_21), .partial_sum_in(reg_psum_50_21), .reg_activation(reg_activation_51_21), .reg_weight(reg_weight_51_21), .reg_partial_sum(reg_psum_51_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_22( .activation_in(reg_activation_51_21), .weight_in(reg_weight_50_22), .partial_sum_in(reg_psum_50_22), .reg_activation(reg_activation_51_22), .reg_weight(reg_weight_51_22), .reg_partial_sum(reg_psum_51_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_23( .activation_in(reg_activation_51_22), .weight_in(reg_weight_50_23), .partial_sum_in(reg_psum_50_23), .reg_activation(reg_activation_51_23), .reg_weight(reg_weight_51_23), .reg_partial_sum(reg_psum_51_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_24( .activation_in(reg_activation_51_23), .weight_in(reg_weight_50_24), .partial_sum_in(reg_psum_50_24), .reg_activation(reg_activation_51_24), .reg_weight(reg_weight_51_24), .reg_partial_sum(reg_psum_51_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_25( .activation_in(reg_activation_51_24), .weight_in(reg_weight_50_25), .partial_sum_in(reg_psum_50_25), .reg_activation(reg_activation_51_25), .reg_weight(reg_weight_51_25), .reg_partial_sum(reg_psum_51_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_26( .activation_in(reg_activation_51_25), .weight_in(reg_weight_50_26), .partial_sum_in(reg_psum_50_26), .reg_activation(reg_activation_51_26), .reg_weight(reg_weight_51_26), .reg_partial_sum(reg_psum_51_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_27( .activation_in(reg_activation_51_26), .weight_in(reg_weight_50_27), .partial_sum_in(reg_psum_50_27), .reg_activation(reg_activation_51_27), .reg_weight(reg_weight_51_27), .reg_partial_sum(reg_psum_51_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_28( .activation_in(reg_activation_51_27), .weight_in(reg_weight_50_28), .partial_sum_in(reg_psum_50_28), .reg_activation(reg_activation_51_28), .reg_weight(reg_weight_51_28), .reg_partial_sum(reg_psum_51_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_29( .activation_in(reg_activation_51_28), .weight_in(reg_weight_50_29), .partial_sum_in(reg_psum_50_29), .reg_activation(reg_activation_51_29), .reg_weight(reg_weight_51_29), .reg_partial_sum(reg_psum_51_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_30( .activation_in(reg_activation_51_29), .weight_in(reg_weight_50_30), .partial_sum_in(reg_psum_50_30), .reg_activation(reg_activation_51_30), .reg_weight(reg_weight_51_30), .reg_partial_sum(reg_psum_51_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_31( .activation_in(reg_activation_51_30), .weight_in(reg_weight_50_31), .partial_sum_in(reg_psum_50_31), .reg_activation(reg_activation_51_31), .reg_weight(reg_weight_51_31), .reg_partial_sum(reg_psum_51_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_32( .activation_in(reg_activation_51_31), .weight_in(reg_weight_50_32), .partial_sum_in(reg_psum_50_32), .reg_activation(reg_activation_51_32), .reg_weight(reg_weight_51_32), .reg_partial_sum(reg_psum_51_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_33( .activation_in(reg_activation_51_32), .weight_in(reg_weight_50_33), .partial_sum_in(reg_psum_50_33), .reg_activation(reg_activation_51_33), .reg_weight(reg_weight_51_33), .reg_partial_sum(reg_psum_51_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_34( .activation_in(reg_activation_51_33), .weight_in(reg_weight_50_34), .partial_sum_in(reg_psum_50_34), .reg_activation(reg_activation_51_34), .reg_weight(reg_weight_51_34), .reg_partial_sum(reg_psum_51_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_35( .activation_in(reg_activation_51_34), .weight_in(reg_weight_50_35), .partial_sum_in(reg_psum_50_35), .reg_activation(reg_activation_51_35), .reg_weight(reg_weight_51_35), .reg_partial_sum(reg_psum_51_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_36( .activation_in(reg_activation_51_35), .weight_in(reg_weight_50_36), .partial_sum_in(reg_psum_50_36), .reg_activation(reg_activation_51_36), .reg_weight(reg_weight_51_36), .reg_partial_sum(reg_psum_51_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_37( .activation_in(reg_activation_51_36), .weight_in(reg_weight_50_37), .partial_sum_in(reg_psum_50_37), .reg_activation(reg_activation_51_37), .reg_weight(reg_weight_51_37), .reg_partial_sum(reg_psum_51_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_38( .activation_in(reg_activation_51_37), .weight_in(reg_weight_50_38), .partial_sum_in(reg_psum_50_38), .reg_activation(reg_activation_51_38), .reg_weight(reg_weight_51_38), .reg_partial_sum(reg_psum_51_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_39( .activation_in(reg_activation_51_38), .weight_in(reg_weight_50_39), .partial_sum_in(reg_psum_50_39), .reg_activation(reg_activation_51_39), .reg_weight(reg_weight_51_39), .reg_partial_sum(reg_psum_51_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_40( .activation_in(reg_activation_51_39), .weight_in(reg_weight_50_40), .partial_sum_in(reg_psum_50_40), .reg_activation(reg_activation_51_40), .reg_weight(reg_weight_51_40), .reg_partial_sum(reg_psum_51_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_41( .activation_in(reg_activation_51_40), .weight_in(reg_weight_50_41), .partial_sum_in(reg_psum_50_41), .reg_activation(reg_activation_51_41), .reg_weight(reg_weight_51_41), .reg_partial_sum(reg_psum_51_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_42( .activation_in(reg_activation_51_41), .weight_in(reg_weight_50_42), .partial_sum_in(reg_psum_50_42), .reg_activation(reg_activation_51_42), .reg_weight(reg_weight_51_42), .reg_partial_sum(reg_psum_51_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_43( .activation_in(reg_activation_51_42), .weight_in(reg_weight_50_43), .partial_sum_in(reg_psum_50_43), .reg_activation(reg_activation_51_43), .reg_weight(reg_weight_51_43), .reg_partial_sum(reg_psum_51_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_44( .activation_in(reg_activation_51_43), .weight_in(reg_weight_50_44), .partial_sum_in(reg_psum_50_44), .reg_activation(reg_activation_51_44), .reg_weight(reg_weight_51_44), .reg_partial_sum(reg_psum_51_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_45( .activation_in(reg_activation_51_44), .weight_in(reg_weight_50_45), .partial_sum_in(reg_psum_50_45), .reg_activation(reg_activation_51_45), .reg_weight(reg_weight_51_45), .reg_partial_sum(reg_psum_51_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_46( .activation_in(reg_activation_51_45), .weight_in(reg_weight_50_46), .partial_sum_in(reg_psum_50_46), .reg_activation(reg_activation_51_46), .reg_weight(reg_weight_51_46), .reg_partial_sum(reg_psum_51_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_47( .activation_in(reg_activation_51_46), .weight_in(reg_weight_50_47), .partial_sum_in(reg_psum_50_47), .reg_activation(reg_activation_51_47), .reg_weight(reg_weight_51_47), .reg_partial_sum(reg_psum_51_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_48( .activation_in(reg_activation_51_47), .weight_in(reg_weight_50_48), .partial_sum_in(reg_psum_50_48), .reg_activation(reg_activation_51_48), .reg_weight(reg_weight_51_48), .reg_partial_sum(reg_psum_51_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_49( .activation_in(reg_activation_51_48), .weight_in(reg_weight_50_49), .partial_sum_in(reg_psum_50_49), .reg_activation(reg_activation_51_49), .reg_weight(reg_weight_51_49), .reg_partial_sum(reg_psum_51_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_50( .activation_in(reg_activation_51_49), .weight_in(reg_weight_50_50), .partial_sum_in(reg_psum_50_50), .reg_activation(reg_activation_51_50), .reg_weight(reg_weight_51_50), .reg_partial_sum(reg_psum_51_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_51( .activation_in(reg_activation_51_50), .weight_in(reg_weight_50_51), .partial_sum_in(reg_psum_50_51), .reg_activation(reg_activation_51_51), .reg_weight(reg_weight_51_51), .reg_partial_sum(reg_psum_51_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_52( .activation_in(reg_activation_51_51), .weight_in(reg_weight_50_52), .partial_sum_in(reg_psum_50_52), .reg_activation(reg_activation_51_52), .reg_weight(reg_weight_51_52), .reg_partial_sum(reg_psum_51_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_53( .activation_in(reg_activation_51_52), .weight_in(reg_weight_50_53), .partial_sum_in(reg_psum_50_53), .reg_activation(reg_activation_51_53), .reg_weight(reg_weight_51_53), .reg_partial_sum(reg_psum_51_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_54( .activation_in(reg_activation_51_53), .weight_in(reg_weight_50_54), .partial_sum_in(reg_psum_50_54), .reg_activation(reg_activation_51_54), .reg_weight(reg_weight_51_54), .reg_partial_sum(reg_psum_51_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_55( .activation_in(reg_activation_51_54), .weight_in(reg_weight_50_55), .partial_sum_in(reg_psum_50_55), .reg_activation(reg_activation_51_55), .reg_weight(reg_weight_51_55), .reg_partial_sum(reg_psum_51_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_56( .activation_in(reg_activation_51_55), .weight_in(reg_weight_50_56), .partial_sum_in(reg_psum_50_56), .reg_activation(reg_activation_51_56), .reg_weight(reg_weight_51_56), .reg_partial_sum(reg_psum_51_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_57( .activation_in(reg_activation_51_56), .weight_in(reg_weight_50_57), .partial_sum_in(reg_psum_50_57), .reg_activation(reg_activation_51_57), .reg_weight(reg_weight_51_57), .reg_partial_sum(reg_psum_51_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_58( .activation_in(reg_activation_51_57), .weight_in(reg_weight_50_58), .partial_sum_in(reg_psum_50_58), .reg_activation(reg_activation_51_58), .reg_weight(reg_weight_51_58), .reg_partial_sum(reg_psum_51_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_59( .activation_in(reg_activation_51_58), .weight_in(reg_weight_50_59), .partial_sum_in(reg_psum_50_59), .reg_activation(reg_activation_51_59), .reg_weight(reg_weight_51_59), .reg_partial_sum(reg_psum_51_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_60( .activation_in(reg_activation_51_59), .weight_in(reg_weight_50_60), .partial_sum_in(reg_psum_50_60), .reg_activation(reg_activation_51_60), .reg_weight(reg_weight_51_60), .reg_partial_sum(reg_psum_51_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_61( .activation_in(reg_activation_51_60), .weight_in(reg_weight_50_61), .partial_sum_in(reg_psum_50_61), .reg_activation(reg_activation_51_61), .reg_weight(reg_weight_51_61), .reg_partial_sum(reg_psum_51_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_62( .activation_in(reg_activation_51_61), .weight_in(reg_weight_50_62), .partial_sum_in(reg_psum_50_62), .reg_activation(reg_activation_51_62), .reg_weight(reg_weight_51_62), .reg_partial_sum(reg_psum_51_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U51_63( .activation_in(reg_activation_51_62), .weight_in(reg_weight_50_63), .partial_sum_in(reg_psum_50_63), .reg_weight(reg_weight_51_63), .reg_partial_sum(reg_psum_51_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_0( .activation_in(in_activation_52), .weight_in(reg_weight_51_0), .partial_sum_in(reg_psum_51_0), .reg_activation(reg_activation_52_0), .reg_weight(reg_weight_52_0), .reg_partial_sum(reg_psum_52_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_1( .activation_in(reg_activation_52_0), .weight_in(reg_weight_51_1), .partial_sum_in(reg_psum_51_1), .reg_activation(reg_activation_52_1), .reg_weight(reg_weight_52_1), .reg_partial_sum(reg_psum_52_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_2( .activation_in(reg_activation_52_1), .weight_in(reg_weight_51_2), .partial_sum_in(reg_psum_51_2), .reg_activation(reg_activation_52_2), .reg_weight(reg_weight_52_2), .reg_partial_sum(reg_psum_52_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_3( .activation_in(reg_activation_52_2), .weight_in(reg_weight_51_3), .partial_sum_in(reg_psum_51_3), .reg_activation(reg_activation_52_3), .reg_weight(reg_weight_52_3), .reg_partial_sum(reg_psum_52_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_4( .activation_in(reg_activation_52_3), .weight_in(reg_weight_51_4), .partial_sum_in(reg_psum_51_4), .reg_activation(reg_activation_52_4), .reg_weight(reg_weight_52_4), .reg_partial_sum(reg_psum_52_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_5( .activation_in(reg_activation_52_4), .weight_in(reg_weight_51_5), .partial_sum_in(reg_psum_51_5), .reg_activation(reg_activation_52_5), .reg_weight(reg_weight_52_5), .reg_partial_sum(reg_psum_52_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_6( .activation_in(reg_activation_52_5), .weight_in(reg_weight_51_6), .partial_sum_in(reg_psum_51_6), .reg_activation(reg_activation_52_6), .reg_weight(reg_weight_52_6), .reg_partial_sum(reg_psum_52_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_7( .activation_in(reg_activation_52_6), .weight_in(reg_weight_51_7), .partial_sum_in(reg_psum_51_7), .reg_activation(reg_activation_52_7), .reg_weight(reg_weight_52_7), .reg_partial_sum(reg_psum_52_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_8( .activation_in(reg_activation_52_7), .weight_in(reg_weight_51_8), .partial_sum_in(reg_psum_51_8), .reg_activation(reg_activation_52_8), .reg_weight(reg_weight_52_8), .reg_partial_sum(reg_psum_52_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_9( .activation_in(reg_activation_52_8), .weight_in(reg_weight_51_9), .partial_sum_in(reg_psum_51_9), .reg_activation(reg_activation_52_9), .reg_weight(reg_weight_52_9), .reg_partial_sum(reg_psum_52_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_10( .activation_in(reg_activation_52_9), .weight_in(reg_weight_51_10), .partial_sum_in(reg_psum_51_10), .reg_activation(reg_activation_52_10), .reg_weight(reg_weight_52_10), .reg_partial_sum(reg_psum_52_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_11( .activation_in(reg_activation_52_10), .weight_in(reg_weight_51_11), .partial_sum_in(reg_psum_51_11), .reg_activation(reg_activation_52_11), .reg_weight(reg_weight_52_11), .reg_partial_sum(reg_psum_52_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_12( .activation_in(reg_activation_52_11), .weight_in(reg_weight_51_12), .partial_sum_in(reg_psum_51_12), .reg_activation(reg_activation_52_12), .reg_weight(reg_weight_52_12), .reg_partial_sum(reg_psum_52_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_13( .activation_in(reg_activation_52_12), .weight_in(reg_weight_51_13), .partial_sum_in(reg_psum_51_13), .reg_activation(reg_activation_52_13), .reg_weight(reg_weight_52_13), .reg_partial_sum(reg_psum_52_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_14( .activation_in(reg_activation_52_13), .weight_in(reg_weight_51_14), .partial_sum_in(reg_psum_51_14), .reg_activation(reg_activation_52_14), .reg_weight(reg_weight_52_14), .reg_partial_sum(reg_psum_52_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_15( .activation_in(reg_activation_52_14), .weight_in(reg_weight_51_15), .partial_sum_in(reg_psum_51_15), .reg_activation(reg_activation_52_15), .reg_weight(reg_weight_52_15), .reg_partial_sum(reg_psum_52_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_16( .activation_in(reg_activation_52_15), .weight_in(reg_weight_51_16), .partial_sum_in(reg_psum_51_16), .reg_activation(reg_activation_52_16), .reg_weight(reg_weight_52_16), .reg_partial_sum(reg_psum_52_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_17( .activation_in(reg_activation_52_16), .weight_in(reg_weight_51_17), .partial_sum_in(reg_psum_51_17), .reg_activation(reg_activation_52_17), .reg_weight(reg_weight_52_17), .reg_partial_sum(reg_psum_52_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_18( .activation_in(reg_activation_52_17), .weight_in(reg_weight_51_18), .partial_sum_in(reg_psum_51_18), .reg_activation(reg_activation_52_18), .reg_weight(reg_weight_52_18), .reg_partial_sum(reg_psum_52_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_19( .activation_in(reg_activation_52_18), .weight_in(reg_weight_51_19), .partial_sum_in(reg_psum_51_19), .reg_activation(reg_activation_52_19), .reg_weight(reg_weight_52_19), .reg_partial_sum(reg_psum_52_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_20( .activation_in(reg_activation_52_19), .weight_in(reg_weight_51_20), .partial_sum_in(reg_psum_51_20), .reg_activation(reg_activation_52_20), .reg_weight(reg_weight_52_20), .reg_partial_sum(reg_psum_52_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_21( .activation_in(reg_activation_52_20), .weight_in(reg_weight_51_21), .partial_sum_in(reg_psum_51_21), .reg_activation(reg_activation_52_21), .reg_weight(reg_weight_52_21), .reg_partial_sum(reg_psum_52_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_22( .activation_in(reg_activation_52_21), .weight_in(reg_weight_51_22), .partial_sum_in(reg_psum_51_22), .reg_activation(reg_activation_52_22), .reg_weight(reg_weight_52_22), .reg_partial_sum(reg_psum_52_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_23( .activation_in(reg_activation_52_22), .weight_in(reg_weight_51_23), .partial_sum_in(reg_psum_51_23), .reg_activation(reg_activation_52_23), .reg_weight(reg_weight_52_23), .reg_partial_sum(reg_psum_52_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_24( .activation_in(reg_activation_52_23), .weight_in(reg_weight_51_24), .partial_sum_in(reg_psum_51_24), .reg_activation(reg_activation_52_24), .reg_weight(reg_weight_52_24), .reg_partial_sum(reg_psum_52_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_25( .activation_in(reg_activation_52_24), .weight_in(reg_weight_51_25), .partial_sum_in(reg_psum_51_25), .reg_activation(reg_activation_52_25), .reg_weight(reg_weight_52_25), .reg_partial_sum(reg_psum_52_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_26( .activation_in(reg_activation_52_25), .weight_in(reg_weight_51_26), .partial_sum_in(reg_psum_51_26), .reg_activation(reg_activation_52_26), .reg_weight(reg_weight_52_26), .reg_partial_sum(reg_psum_52_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_27( .activation_in(reg_activation_52_26), .weight_in(reg_weight_51_27), .partial_sum_in(reg_psum_51_27), .reg_activation(reg_activation_52_27), .reg_weight(reg_weight_52_27), .reg_partial_sum(reg_psum_52_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_28( .activation_in(reg_activation_52_27), .weight_in(reg_weight_51_28), .partial_sum_in(reg_psum_51_28), .reg_activation(reg_activation_52_28), .reg_weight(reg_weight_52_28), .reg_partial_sum(reg_psum_52_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_29( .activation_in(reg_activation_52_28), .weight_in(reg_weight_51_29), .partial_sum_in(reg_psum_51_29), .reg_activation(reg_activation_52_29), .reg_weight(reg_weight_52_29), .reg_partial_sum(reg_psum_52_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_30( .activation_in(reg_activation_52_29), .weight_in(reg_weight_51_30), .partial_sum_in(reg_psum_51_30), .reg_activation(reg_activation_52_30), .reg_weight(reg_weight_52_30), .reg_partial_sum(reg_psum_52_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_31( .activation_in(reg_activation_52_30), .weight_in(reg_weight_51_31), .partial_sum_in(reg_psum_51_31), .reg_activation(reg_activation_52_31), .reg_weight(reg_weight_52_31), .reg_partial_sum(reg_psum_52_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_32( .activation_in(reg_activation_52_31), .weight_in(reg_weight_51_32), .partial_sum_in(reg_psum_51_32), .reg_activation(reg_activation_52_32), .reg_weight(reg_weight_52_32), .reg_partial_sum(reg_psum_52_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_33( .activation_in(reg_activation_52_32), .weight_in(reg_weight_51_33), .partial_sum_in(reg_psum_51_33), .reg_activation(reg_activation_52_33), .reg_weight(reg_weight_52_33), .reg_partial_sum(reg_psum_52_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_34( .activation_in(reg_activation_52_33), .weight_in(reg_weight_51_34), .partial_sum_in(reg_psum_51_34), .reg_activation(reg_activation_52_34), .reg_weight(reg_weight_52_34), .reg_partial_sum(reg_psum_52_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_35( .activation_in(reg_activation_52_34), .weight_in(reg_weight_51_35), .partial_sum_in(reg_psum_51_35), .reg_activation(reg_activation_52_35), .reg_weight(reg_weight_52_35), .reg_partial_sum(reg_psum_52_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_36( .activation_in(reg_activation_52_35), .weight_in(reg_weight_51_36), .partial_sum_in(reg_psum_51_36), .reg_activation(reg_activation_52_36), .reg_weight(reg_weight_52_36), .reg_partial_sum(reg_psum_52_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_37( .activation_in(reg_activation_52_36), .weight_in(reg_weight_51_37), .partial_sum_in(reg_psum_51_37), .reg_activation(reg_activation_52_37), .reg_weight(reg_weight_52_37), .reg_partial_sum(reg_psum_52_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_38( .activation_in(reg_activation_52_37), .weight_in(reg_weight_51_38), .partial_sum_in(reg_psum_51_38), .reg_activation(reg_activation_52_38), .reg_weight(reg_weight_52_38), .reg_partial_sum(reg_psum_52_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_39( .activation_in(reg_activation_52_38), .weight_in(reg_weight_51_39), .partial_sum_in(reg_psum_51_39), .reg_activation(reg_activation_52_39), .reg_weight(reg_weight_52_39), .reg_partial_sum(reg_psum_52_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_40( .activation_in(reg_activation_52_39), .weight_in(reg_weight_51_40), .partial_sum_in(reg_psum_51_40), .reg_activation(reg_activation_52_40), .reg_weight(reg_weight_52_40), .reg_partial_sum(reg_psum_52_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_41( .activation_in(reg_activation_52_40), .weight_in(reg_weight_51_41), .partial_sum_in(reg_psum_51_41), .reg_activation(reg_activation_52_41), .reg_weight(reg_weight_52_41), .reg_partial_sum(reg_psum_52_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_42( .activation_in(reg_activation_52_41), .weight_in(reg_weight_51_42), .partial_sum_in(reg_psum_51_42), .reg_activation(reg_activation_52_42), .reg_weight(reg_weight_52_42), .reg_partial_sum(reg_psum_52_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_43( .activation_in(reg_activation_52_42), .weight_in(reg_weight_51_43), .partial_sum_in(reg_psum_51_43), .reg_activation(reg_activation_52_43), .reg_weight(reg_weight_52_43), .reg_partial_sum(reg_psum_52_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_44( .activation_in(reg_activation_52_43), .weight_in(reg_weight_51_44), .partial_sum_in(reg_psum_51_44), .reg_activation(reg_activation_52_44), .reg_weight(reg_weight_52_44), .reg_partial_sum(reg_psum_52_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_45( .activation_in(reg_activation_52_44), .weight_in(reg_weight_51_45), .partial_sum_in(reg_psum_51_45), .reg_activation(reg_activation_52_45), .reg_weight(reg_weight_52_45), .reg_partial_sum(reg_psum_52_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_46( .activation_in(reg_activation_52_45), .weight_in(reg_weight_51_46), .partial_sum_in(reg_psum_51_46), .reg_activation(reg_activation_52_46), .reg_weight(reg_weight_52_46), .reg_partial_sum(reg_psum_52_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_47( .activation_in(reg_activation_52_46), .weight_in(reg_weight_51_47), .partial_sum_in(reg_psum_51_47), .reg_activation(reg_activation_52_47), .reg_weight(reg_weight_52_47), .reg_partial_sum(reg_psum_52_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_48( .activation_in(reg_activation_52_47), .weight_in(reg_weight_51_48), .partial_sum_in(reg_psum_51_48), .reg_activation(reg_activation_52_48), .reg_weight(reg_weight_52_48), .reg_partial_sum(reg_psum_52_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_49( .activation_in(reg_activation_52_48), .weight_in(reg_weight_51_49), .partial_sum_in(reg_psum_51_49), .reg_activation(reg_activation_52_49), .reg_weight(reg_weight_52_49), .reg_partial_sum(reg_psum_52_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_50( .activation_in(reg_activation_52_49), .weight_in(reg_weight_51_50), .partial_sum_in(reg_psum_51_50), .reg_activation(reg_activation_52_50), .reg_weight(reg_weight_52_50), .reg_partial_sum(reg_psum_52_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_51( .activation_in(reg_activation_52_50), .weight_in(reg_weight_51_51), .partial_sum_in(reg_psum_51_51), .reg_activation(reg_activation_52_51), .reg_weight(reg_weight_52_51), .reg_partial_sum(reg_psum_52_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_52( .activation_in(reg_activation_52_51), .weight_in(reg_weight_51_52), .partial_sum_in(reg_psum_51_52), .reg_activation(reg_activation_52_52), .reg_weight(reg_weight_52_52), .reg_partial_sum(reg_psum_52_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_53( .activation_in(reg_activation_52_52), .weight_in(reg_weight_51_53), .partial_sum_in(reg_psum_51_53), .reg_activation(reg_activation_52_53), .reg_weight(reg_weight_52_53), .reg_partial_sum(reg_psum_52_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_54( .activation_in(reg_activation_52_53), .weight_in(reg_weight_51_54), .partial_sum_in(reg_psum_51_54), .reg_activation(reg_activation_52_54), .reg_weight(reg_weight_52_54), .reg_partial_sum(reg_psum_52_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_55( .activation_in(reg_activation_52_54), .weight_in(reg_weight_51_55), .partial_sum_in(reg_psum_51_55), .reg_activation(reg_activation_52_55), .reg_weight(reg_weight_52_55), .reg_partial_sum(reg_psum_52_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_56( .activation_in(reg_activation_52_55), .weight_in(reg_weight_51_56), .partial_sum_in(reg_psum_51_56), .reg_activation(reg_activation_52_56), .reg_weight(reg_weight_52_56), .reg_partial_sum(reg_psum_52_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_57( .activation_in(reg_activation_52_56), .weight_in(reg_weight_51_57), .partial_sum_in(reg_psum_51_57), .reg_activation(reg_activation_52_57), .reg_weight(reg_weight_52_57), .reg_partial_sum(reg_psum_52_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_58( .activation_in(reg_activation_52_57), .weight_in(reg_weight_51_58), .partial_sum_in(reg_psum_51_58), .reg_activation(reg_activation_52_58), .reg_weight(reg_weight_52_58), .reg_partial_sum(reg_psum_52_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_59( .activation_in(reg_activation_52_58), .weight_in(reg_weight_51_59), .partial_sum_in(reg_psum_51_59), .reg_activation(reg_activation_52_59), .reg_weight(reg_weight_52_59), .reg_partial_sum(reg_psum_52_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_60( .activation_in(reg_activation_52_59), .weight_in(reg_weight_51_60), .partial_sum_in(reg_psum_51_60), .reg_activation(reg_activation_52_60), .reg_weight(reg_weight_52_60), .reg_partial_sum(reg_psum_52_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_61( .activation_in(reg_activation_52_60), .weight_in(reg_weight_51_61), .partial_sum_in(reg_psum_51_61), .reg_activation(reg_activation_52_61), .reg_weight(reg_weight_52_61), .reg_partial_sum(reg_psum_52_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_62( .activation_in(reg_activation_52_61), .weight_in(reg_weight_51_62), .partial_sum_in(reg_psum_51_62), .reg_activation(reg_activation_52_62), .reg_weight(reg_weight_52_62), .reg_partial_sum(reg_psum_52_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U52_63( .activation_in(reg_activation_52_62), .weight_in(reg_weight_51_63), .partial_sum_in(reg_psum_51_63), .reg_weight(reg_weight_52_63), .reg_partial_sum(reg_psum_52_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_0( .activation_in(in_activation_53), .weight_in(reg_weight_52_0), .partial_sum_in(reg_psum_52_0), .reg_activation(reg_activation_53_0), .reg_weight(reg_weight_53_0), .reg_partial_sum(reg_psum_53_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_1( .activation_in(reg_activation_53_0), .weight_in(reg_weight_52_1), .partial_sum_in(reg_psum_52_1), .reg_activation(reg_activation_53_1), .reg_weight(reg_weight_53_1), .reg_partial_sum(reg_psum_53_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_2( .activation_in(reg_activation_53_1), .weight_in(reg_weight_52_2), .partial_sum_in(reg_psum_52_2), .reg_activation(reg_activation_53_2), .reg_weight(reg_weight_53_2), .reg_partial_sum(reg_psum_53_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_3( .activation_in(reg_activation_53_2), .weight_in(reg_weight_52_3), .partial_sum_in(reg_psum_52_3), .reg_activation(reg_activation_53_3), .reg_weight(reg_weight_53_3), .reg_partial_sum(reg_psum_53_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_4( .activation_in(reg_activation_53_3), .weight_in(reg_weight_52_4), .partial_sum_in(reg_psum_52_4), .reg_activation(reg_activation_53_4), .reg_weight(reg_weight_53_4), .reg_partial_sum(reg_psum_53_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_5( .activation_in(reg_activation_53_4), .weight_in(reg_weight_52_5), .partial_sum_in(reg_psum_52_5), .reg_activation(reg_activation_53_5), .reg_weight(reg_weight_53_5), .reg_partial_sum(reg_psum_53_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_6( .activation_in(reg_activation_53_5), .weight_in(reg_weight_52_6), .partial_sum_in(reg_psum_52_6), .reg_activation(reg_activation_53_6), .reg_weight(reg_weight_53_6), .reg_partial_sum(reg_psum_53_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_7( .activation_in(reg_activation_53_6), .weight_in(reg_weight_52_7), .partial_sum_in(reg_psum_52_7), .reg_activation(reg_activation_53_7), .reg_weight(reg_weight_53_7), .reg_partial_sum(reg_psum_53_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_8( .activation_in(reg_activation_53_7), .weight_in(reg_weight_52_8), .partial_sum_in(reg_psum_52_8), .reg_activation(reg_activation_53_8), .reg_weight(reg_weight_53_8), .reg_partial_sum(reg_psum_53_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_9( .activation_in(reg_activation_53_8), .weight_in(reg_weight_52_9), .partial_sum_in(reg_psum_52_9), .reg_activation(reg_activation_53_9), .reg_weight(reg_weight_53_9), .reg_partial_sum(reg_psum_53_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_10( .activation_in(reg_activation_53_9), .weight_in(reg_weight_52_10), .partial_sum_in(reg_psum_52_10), .reg_activation(reg_activation_53_10), .reg_weight(reg_weight_53_10), .reg_partial_sum(reg_psum_53_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_11( .activation_in(reg_activation_53_10), .weight_in(reg_weight_52_11), .partial_sum_in(reg_psum_52_11), .reg_activation(reg_activation_53_11), .reg_weight(reg_weight_53_11), .reg_partial_sum(reg_psum_53_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_12( .activation_in(reg_activation_53_11), .weight_in(reg_weight_52_12), .partial_sum_in(reg_psum_52_12), .reg_activation(reg_activation_53_12), .reg_weight(reg_weight_53_12), .reg_partial_sum(reg_psum_53_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_13( .activation_in(reg_activation_53_12), .weight_in(reg_weight_52_13), .partial_sum_in(reg_psum_52_13), .reg_activation(reg_activation_53_13), .reg_weight(reg_weight_53_13), .reg_partial_sum(reg_psum_53_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_14( .activation_in(reg_activation_53_13), .weight_in(reg_weight_52_14), .partial_sum_in(reg_psum_52_14), .reg_activation(reg_activation_53_14), .reg_weight(reg_weight_53_14), .reg_partial_sum(reg_psum_53_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_15( .activation_in(reg_activation_53_14), .weight_in(reg_weight_52_15), .partial_sum_in(reg_psum_52_15), .reg_activation(reg_activation_53_15), .reg_weight(reg_weight_53_15), .reg_partial_sum(reg_psum_53_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_16( .activation_in(reg_activation_53_15), .weight_in(reg_weight_52_16), .partial_sum_in(reg_psum_52_16), .reg_activation(reg_activation_53_16), .reg_weight(reg_weight_53_16), .reg_partial_sum(reg_psum_53_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_17( .activation_in(reg_activation_53_16), .weight_in(reg_weight_52_17), .partial_sum_in(reg_psum_52_17), .reg_activation(reg_activation_53_17), .reg_weight(reg_weight_53_17), .reg_partial_sum(reg_psum_53_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_18( .activation_in(reg_activation_53_17), .weight_in(reg_weight_52_18), .partial_sum_in(reg_psum_52_18), .reg_activation(reg_activation_53_18), .reg_weight(reg_weight_53_18), .reg_partial_sum(reg_psum_53_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_19( .activation_in(reg_activation_53_18), .weight_in(reg_weight_52_19), .partial_sum_in(reg_psum_52_19), .reg_activation(reg_activation_53_19), .reg_weight(reg_weight_53_19), .reg_partial_sum(reg_psum_53_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_20( .activation_in(reg_activation_53_19), .weight_in(reg_weight_52_20), .partial_sum_in(reg_psum_52_20), .reg_activation(reg_activation_53_20), .reg_weight(reg_weight_53_20), .reg_partial_sum(reg_psum_53_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_21( .activation_in(reg_activation_53_20), .weight_in(reg_weight_52_21), .partial_sum_in(reg_psum_52_21), .reg_activation(reg_activation_53_21), .reg_weight(reg_weight_53_21), .reg_partial_sum(reg_psum_53_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_22( .activation_in(reg_activation_53_21), .weight_in(reg_weight_52_22), .partial_sum_in(reg_psum_52_22), .reg_activation(reg_activation_53_22), .reg_weight(reg_weight_53_22), .reg_partial_sum(reg_psum_53_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_23( .activation_in(reg_activation_53_22), .weight_in(reg_weight_52_23), .partial_sum_in(reg_psum_52_23), .reg_activation(reg_activation_53_23), .reg_weight(reg_weight_53_23), .reg_partial_sum(reg_psum_53_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_24( .activation_in(reg_activation_53_23), .weight_in(reg_weight_52_24), .partial_sum_in(reg_psum_52_24), .reg_activation(reg_activation_53_24), .reg_weight(reg_weight_53_24), .reg_partial_sum(reg_psum_53_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_25( .activation_in(reg_activation_53_24), .weight_in(reg_weight_52_25), .partial_sum_in(reg_psum_52_25), .reg_activation(reg_activation_53_25), .reg_weight(reg_weight_53_25), .reg_partial_sum(reg_psum_53_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_26( .activation_in(reg_activation_53_25), .weight_in(reg_weight_52_26), .partial_sum_in(reg_psum_52_26), .reg_activation(reg_activation_53_26), .reg_weight(reg_weight_53_26), .reg_partial_sum(reg_psum_53_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_27( .activation_in(reg_activation_53_26), .weight_in(reg_weight_52_27), .partial_sum_in(reg_psum_52_27), .reg_activation(reg_activation_53_27), .reg_weight(reg_weight_53_27), .reg_partial_sum(reg_psum_53_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_28( .activation_in(reg_activation_53_27), .weight_in(reg_weight_52_28), .partial_sum_in(reg_psum_52_28), .reg_activation(reg_activation_53_28), .reg_weight(reg_weight_53_28), .reg_partial_sum(reg_psum_53_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_29( .activation_in(reg_activation_53_28), .weight_in(reg_weight_52_29), .partial_sum_in(reg_psum_52_29), .reg_activation(reg_activation_53_29), .reg_weight(reg_weight_53_29), .reg_partial_sum(reg_psum_53_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_30( .activation_in(reg_activation_53_29), .weight_in(reg_weight_52_30), .partial_sum_in(reg_psum_52_30), .reg_activation(reg_activation_53_30), .reg_weight(reg_weight_53_30), .reg_partial_sum(reg_psum_53_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_31( .activation_in(reg_activation_53_30), .weight_in(reg_weight_52_31), .partial_sum_in(reg_psum_52_31), .reg_activation(reg_activation_53_31), .reg_weight(reg_weight_53_31), .reg_partial_sum(reg_psum_53_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_32( .activation_in(reg_activation_53_31), .weight_in(reg_weight_52_32), .partial_sum_in(reg_psum_52_32), .reg_activation(reg_activation_53_32), .reg_weight(reg_weight_53_32), .reg_partial_sum(reg_psum_53_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_33( .activation_in(reg_activation_53_32), .weight_in(reg_weight_52_33), .partial_sum_in(reg_psum_52_33), .reg_activation(reg_activation_53_33), .reg_weight(reg_weight_53_33), .reg_partial_sum(reg_psum_53_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_34( .activation_in(reg_activation_53_33), .weight_in(reg_weight_52_34), .partial_sum_in(reg_psum_52_34), .reg_activation(reg_activation_53_34), .reg_weight(reg_weight_53_34), .reg_partial_sum(reg_psum_53_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_35( .activation_in(reg_activation_53_34), .weight_in(reg_weight_52_35), .partial_sum_in(reg_psum_52_35), .reg_activation(reg_activation_53_35), .reg_weight(reg_weight_53_35), .reg_partial_sum(reg_psum_53_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_36( .activation_in(reg_activation_53_35), .weight_in(reg_weight_52_36), .partial_sum_in(reg_psum_52_36), .reg_activation(reg_activation_53_36), .reg_weight(reg_weight_53_36), .reg_partial_sum(reg_psum_53_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_37( .activation_in(reg_activation_53_36), .weight_in(reg_weight_52_37), .partial_sum_in(reg_psum_52_37), .reg_activation(reg_activation_53_37), .reg_weight(reg_weight_53_37), .reg_partial_sum(reg_psum_53_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_38( .activation_in(reg_activation_53_37), .weight_in(reg_weight_52_38), .partial_sum_in(reg_psum_52_38), .reg_activation(reg_activation_53_38), .reg_weight(reg_weight_53_38), .reg_partial_sum(reg_psum_53_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_39( .activation_in(reg_activation_53_38), .weight_in(reg_weight_52_39), .partial_sum_in(reg_psum_52_39), .reg_activation(reg_activation_53_39), .reg_weight(reg_weight_53_39), .reg_partial_sum(reg_psum_53_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_40( .activation_in(reg_activation_53_39), .weight_in(reg_weight_52_40), .partial_sum_in(reg_psum_52_40), .reg_activation(reg_activation_53_40), .reg_weight(reg_weight_53_40), .reg_partial_sum(reg_psum_53_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_41( .activation_in(reg_activation_53_40), .weight_in(reg_weight_52_41), .partial_sum_in(reg_psum_52_41), .reg_activation(reg_activation_53_41), .reg_weight(reg_weight_53_41), .reg_partial_sum(reg_psum_53_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_42( .activation_in(reg_activation_53_41), .weight_in(reg_weight_52_42), .partial_sum_in(reg_psum_52_42), .reg_activation(reg_activation_53_42), .reg_weight(reg_weight_53_42), .reg_partial_sum(reg_psum_53_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_43( .activation_in(reg_activation_53_42), .weight_in(reg_weight_52_43), .partial_sum_in(reg_psum_52_43), .reg_activation(reg_activation_53_43), .reg_weight(reg_weight_53_43), .reg_partial_sum(reg_psum_53_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_44( .activation_in(reg_activation_53_43), .weight_in(reg_weight_52_44), .partial_sum_in(reg_psum_52_44), .reg_activation(reg_activation_53_44), .reg_weight(reg_weight_53_44), .reg_partial_sum(reg_psum_53_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_45( .activation_in(reg_activation_53_44), .weight_in(reg_weight_52_45), .partial_sum_in(reg_psum_52_45), .reg_activation(reg_activation_53_45), .reg_weight(reg_weight_53_45), .reg_partial_sum(reg_psum_53_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_46( .activation_in(reg_activation_53_45), .weight_in(reg_weight_52_46), .partial_sum_in(reg_psum_52_46), .reg_activation(reg_activation_53_46), .reg_weight(reg_weight_53_46), .reg_partial_sum(reg_psum_53_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_47( .activation_in(reg_activation_53_46), .weight_in(reg_weight_52_47), .partial_sum_in(reg_psum_52_47), .reg_activation(reg_activation_53_47), .reg_weight(reg_weight_53_47), .reg_partial_sum(reg_psum_53_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_48( .activation_in(reg_activation_53_47), .weight_in(reg_weight_52_48), .partial_sum_in(reg_psum_52_48), .reg_activation(reg_activation_53_48), .reg_weight(reg_weight_53_48), .reg_partial_sum(reg_psum_53_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_49( .activation_in(reg_activation_53_48), .weight_in(reg_weight_52_49), .partial_sum_in(reg_psum_52_49), .reg_activation(reg_activation_53_49), .reg_weight(reg_weight_53_49), .reg_partial_sum(reg_psum_53_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_50( .activation_in(reg_activation_53_49), .weight_in(reg_weight_52_50), .partial_sum_in(reg_psum_52_50), .reg_activation(reg_activation_53_50), .reg_weight(reg_weight_53_50), .reg_partial_sum(reg_psum_53_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_51( .activation_in(reg_activation_53_50), .weight_in(reg_weight_52_51), .partial_sum_in(reg_psum_52_51), .reg_activation(reg_activation_53_51), .reg_weight(reg_weight_53_51), .reg_partial_sum(reg_psum_53_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_52( .activation_in(reg_activation_53_51), .weight_in(reg_weight_52_52), .partial_sum_in(reg_psum_52_52), .reg_activation(reg_activation_53_52), .reg_weight(reg_weight_53_52), .reg_partial_sum(reg_psum_53_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_53( .activation_in(reg_activation_53_52), .weight_in(reg_weight_52_53), .partial_sum_in(reg_psum_52_53), .reg_activation(reg_activation_53_53), .reg_weight(reg_weight_53_53), .reg_partial_sum(reg_psum_53_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_54( .activation_in(reg_activation_53_53), .weight_in(reg_weight_52_54), .partial_sum_in(reg_psum_52_54), .reg_activation(reg_activation_53_54), .reg_weight(reg_weight_53_54), .reg_partial_sum(reg_psum_53_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_55( .activation_in(reg_activation_53_54), .weight_in(reg_weight_52_55), .partial_sum_in(reg_psum_52_55), .reg_activation(reg_activation_53_55), .reg_weight(reg_weight_53_55), .reg_partial_sum(reg_psum_53_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_56( .activation_in(reg_activation_53_55), .weight_in(reg_weight_52_56), .partial_sum_in(reg_psum_52_56), .reg_activation(reg_activation_53_56), .reg_weight(reg_weight_53_56), .reg_partial_sum(reg_psum_53_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_57( .activation_in(reg_activation_53_56), .weight_in(reg_weight_52_57), .partial_sum_in(reg_psum_52_57), .reg_activation(reg_activation_53_57), .reg_weight(reg_weight_53_57), .reg_partial_sum(reg_psum_53_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_58( .activation_in(reg_activation_53_57), .weight_in(reg_weight_52_58), .partial_sum_in(reg_psum_52_58), .reg_activation(reg_activation_53_58), .reg_weight(reg_weight_53_58), .reg_partial_sum(reg_psum_53_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_59( .activation_in(reg_activation_53_58), .weight_in(reg_weight_52_59), .partial_sum_in(reg_psum_52_59), .reg_activation(reg_activation_53_59), .reg_weight(reg_weight_53_59), .reg_partial_sum(reg_psum_53_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_60( .activation_in(reg_activation_53_59), .weight_in(reg_weight_52_60), .partial_sum_in(reg_psum_52_60), .reg_activation(reg_activation_53_60), .reg_weight(reg_weight_53_60), .reg_partial_sum(reg_psum_53_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_61( .activation_in(reg_activation_53_60), .weight_in(reg_weight_52_61), .partial_sum_in(reg_psum_52_61), .reg_activation(reg_activation_53_61), .reg_weight(reg_weight_53_61), .reg_partial_sum(reg_psum_53_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_62( .activation_in(reg_activation_53_61), .weight_in(reg_weight_52_62), .partial_sum_in(reg_psum_52_62), .reg_activation(reg_activation_53_62), .reg_weight(reg_weight_53_62), .reg_partial_sum(reg_psum_53_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U53_63( .activation_in(reg_activation_53_62), .weight_in(reg_weight_52_63), .partial_sum_in(reg_psum_52_63), .reg_weight(reg_weight_53_63), .reg_partial_sum(reg_psum_53_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_0( .activation_in(in_activation_54), .weight_in(reg_weight_53_0), .partial_sum_in(reg_psum_53_0), .reg_activation(reg_activation_54_0), .reg_weight(reg_weight_54_0), .reg_partial_sum(reg_psum_54_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_1( .activation_in(reg_activation_54_0), .weight_in(reg_weight_53_1), .partial_sum_in(reg_psum_53_1), .reg_activation(reg_activation_54_1), .reg_weight(reg_weight_54_1), .reg_partial_sum(reg_psum_54_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_2( .activation_in(reg_activation_54_1), .weight_in(reg_weight_53_2), .partial_sum_in(reg_psum_53_2), .reg_activation(reg_activation_54_2), .reg_weight(reg_weight_54_2), .reg_partial_sum(reg_psum_54_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_3( .activation_in(reg_activation_54_2), .weight_in(reg_weight_53_3), .partial_sum_in(reg_psum_53_3), .reg_activation(reg_activation_54_3), .reg_weight(reg_weight_54_3), .reg_partial_sum(reg_psum_54_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_4( .activation_in(reg_activation_54_3), .weight_in(reg_weight_53_4), .partial_sum_in(reg_psum_53_4), .reg_activation(reg_activation_54_4), .reg_weight(reg_weight_54_4), .reg_partial_sum(reg_psum_54_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_5( .activation_in(reg_activation_54_4), .weight_in(reg_weight_53_5), .partial_sum_in(reg_psum_53_5), .reg_activation(reg_activation_54_5), .reg_weight(reg_weight_54_5), .reg_partial_sum(reg_psum_54_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_6( .activation_in(reg_activation_54_5), .weight_in(reg_weight_53_6), .partial_sum_in(reg_psum_53_6), .reg_activation(reg_activation_54_6), .reg_weight(reg_weight_54_6), .reg_partial_sum(reg_psum_54_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_7( .activation_in(reg_activation_54_6), .weight_in(reg_weight_53_7), .partial_sum_in(reg_psum_53_7), .reg_activation(reg_activation_54_7), .reg_weight(reg_weight_54_7), .reg_partial_sum(reg_psum_54_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_8( .activation_in(reg_activation_54_7), .weight_in(reg_weight_53_8), .partial_sum_in(reg_psum_53_8), .reg_activation(reg_activation_54_8), .reg_weight(reg_weight_54_8), .reg_partial_sum(reg_psum_54_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_9( .activation_in(reg_activation_54_8), .weight_in(reg_weight_53_9), .partial_sum_in(reg_psum_53_9), .reg_activation(reg_activation_54_9), .reg_weight(reg_weight_54_9), .reg_partial_sum(reg_psum_54_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_10( .activation_in(reg_activation_54_9), .weight_in(reg_weight_53_10), .partial_sum_in(reg_psum_53_10), .reg_activation(reg_activation_54_10), .reg_weight(reg_weight_54_10), .reg_partial_sum(reg_psum_54_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_11( .activation_in(reg_activation_54_10), .weight_in(reg_weight_53_11), .partial_sum_in(reg_psum_53_11), .reg_activation(reg_activation_54_11), .reg_weight(reg_weight_54_11), .reg_partial_sum(reg_psum_54_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_12( .activation_in(reg_activation_54_11), .weight_in(reg_weight_53_12), .partial_sum_in(reg_psum_53_12), .reg_activation(reg_activation_54_12), .reg_weight(reg_weight_54_12), .reg_partial_sum(reg_psum_54_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_13( .activation_in(reg_activation_54_12), .weight_in(reg_weight_53_13), .partial_sum_in(reg_psum_53_13), .reg_activation(reg_activation_54_13), .reg_weight(reg_weight_54_13), .reg_partial_sum(reg_psum_54_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_14( .activation_in(reg_activation_54_13), .weight_in(reg_weight_53_14), .partial_sum_in(reg_psum_53_14), .reg_activation(reg_activation_54_14), .reg_weight(reg_weight_54_14), .reg_partial_sum(reg_psum_54_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_15( .activation_in(reg_activation_54_14), .weight_in(reg_weight_53_15), .partial_sum_in(reg_psum_53_15), .reg_activation(reg_activation_54_15), .reg_weight(reg_weight_54_15), .reg_partial_sum(reg_psum_54_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_16( .activation_in(reg_activation_54_15), .weight_in(reg_weight_53_16), .partial_sum_in(reg_psum_53_16), .reg_activation(reg_activation_54_16), .reg_weight(reg_weight_54_16), .reg_partial_sum(reg_psum_54_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_17( .activation_in(reg_activation_54_16), .weight_in(reg_weight_53_17), .partial_sum_in(reg_psum_53_17), .reg_activation(reg_activation_54_17), .reg_weight(reg_weight_54_17), .reg_partial_sum(reg_psum_54_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_18( .activation_in(reg_activation_54_17), .weight_in(reg_weight_53_18), .partial_sum_in(reg_psum_53_18), .reg_activation(reg_activation_54_18), .reg_weight(reg_weight_54_18), .reg_partial_sum(reg_psum_54_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_19( .activation_in(reg_activation_54_18), .weight_in(reg_weight_53_19), .partial_sum_in(reg_psum_53_19), .reg_activation(reg_activation_54_19), .reg_weight(reg_weight_54_19), .reg_partial_sum(reg_psum_54_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_20( .activation_in(reg_activation_54_19), .weight_in(reg_weight_53_20), .partial_sum_in(reg_psum_53_20), .reg_activation(reg_activation_54_20), .reg_weight(reg_weight_54_20), .reg_partial_sum(reg_psum_54_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_21( .activation_in(reg_activation_54_20), .weight_in(reg_weight_53_21), .partial_sum_in(reg_psum_53_21), .reg_activation(reg_activation_54_21), .reg_weight(reg_weight_54_21), .reg_partial_sum(reg_psum_54_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_22( .activation_in(reg_activation_54_21), .weight_in(reg_weight_53_22), .partial_sum_in(reg_psum_53_22), .reg_activation(reg_activation_54_22), .reg_weight(reg_weight_54_22), .reg_partial_sum(reg_psum_54_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_23( .activation_in(reg_activation_54_22), .weight_in(reg_weight_53_23), .partial_sum_in(reg_psum_53_23), .reg_activation(reg_activation_54_23), .reg_weight(reg_weight_54_23), .reg_partial_sum(reg_psum_54_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_24( .activation_in(reg_activation_54_23), .weight_in(reg_weight_53_24), .partial_sum_in(reg_psum_53_24), .reg_activation(reg_activation_54_24), .reg_weight(reg_weight_54_24), .reg_partial_sum(reg_psum_54_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_25( .activation_in(reg_activation_54_24), .weight_in(reg_weight_53_25), .partial_sum_in(reg_psum_53_25), .reg_activation(reg_activation_54_25), .reg_weight(reg_weight_54_25), .reg_partial_sum(reg_psum_54_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_26( .activation_in(reg_activation_54_25), .weight_in(reg_weight_53_26), .partial_sum_in(reg_psum_53_26), .reg_activation(reg_activation_54_26), .reg_weight(reg_weight_54_26), .reg_partial_sum(reg_psum_54_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_27( .activation_in(reg_activation_54_26), .weight_in(reg_weight_53_27), .partial_sum_in(reg_psum_53_27), .reg_activation(reg_activation_54_27), .reg_weight(reg_weight_54_27), .reg_partial_sum(reg_psum_54_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_28( .activation_in(reg_activation_54_27), .weight_in(reg_weight_53_28), .partial_sum_in(reg_psum_53_28), .reg_activation(reg_activation_54_28), .reg_weight(reg_weight_54_28), .reg_partial_sum(reg_psum_54_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_29( .activation_in(reg_activation_54_28), .weight_in(reg_weight_53_29), .partial_sum_in(reg_psum_53_29), .reg_activation(reg_activation_54_29), .reg_weight(reg_weight_54_29), .reg_partial_sum(reg_psum_54_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_30( .activation_in(reg_activation_54_29), .weight_in(reg_weight_53_30), .partial_sum_in(reg_psum_53_30), .reg_activation(reg_activation_54_30), .reg_weight(reg_weight_54_30), .reg_partial_sum(reg_psum_54_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_31( .activation_in(reg_activation_54_30), .weight_in(reg_weight_53_31), .partial_sum_in(reg_psum_53_31), .reg_activation(reg_activation_54_31), .reg_weight(reg_weight_54_31), .reg_partial_sum(reg_psum_54_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_32( .activation_in(reg_activation_54_31), .weight_in(reg_weight_53_32), .partial_sum_in(reg_psum_53_32), .reg_activation(reg_activation_54_32), .reg_weight(reg_weight_54_32), .reg_partial_sum(reg_psum_54_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_33( .activation_in(reg_activation_54_32), .weight_in(reg_weight_53_33), .partial_sum_in(reg_psum_53_33), .reg_activation(reg_activation_54_33), .reg_weight(reg_weight_54_33), .reg_partial_sum(reg_psum_54_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_34( .activation_in(reg_activation_54_33), .weight_in(reg_weight_53_34), .partial_sum_in(reg_psum_53_34), .reg_activation(reg_activation_54_34), .reg_weight(reg_weight_54_34), .reg_partial_sum(reg_psum_54_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_35( .activation_in(reg_activation_54_34), .weight_in(reg_weight_53_35), .partial_sum_in(reg_psum_53_35), .reg_activation(reg_activation_54_35), .reg_weight(reg_weight_54_35), .reg_partial_sum(reg_psum_54_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_36( .activation_in(reg_activation_54_35), .weight_in(reg_weight_53_36), .partial_sum_in(reg_psum_53_36), .reg_activation(reg_activation_54_36), .reg_weight(reg_weight_54_36), .reg_partial_sum(reg_psum_54_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_37( .activation_in(reg_activation_54_36), .weight_in(reg_weight_53_37), .partial_sum_in(reg_psum_53_37), .reg_activation(reg_activation_54_37), .reg_weight(reg_weight_54_37), .reg_partial_sum(reg_psum_54_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_38( .activation_in(reg_activation_54_37), .weight_in(reg_weight_53_38), .partial_sum_in(reg_psum_53_38), .reg_activation(reg_activation_54_38), .reg_weight(reg_weight_54_38), .reg_partial_sum(reg_psum_54_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_39( .activation_in(reg_activation_54_38), .weight_in(reg_weight_53_39), .partial_sum_in(reg_psum_53_39), .reg_activation(reg_activation_54_39), .reg_weight(reg_weight_54_39), .reg_partial_sum(reg_psum_54_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_40( .activation_in(reg_activation_54_39), .weight_in(reg_weight_53_40), .partial_sum_in(reg_psum_53_40), .reg_activation(reg_activation_54_40), .reg_weight(reg_weight_54_40), .reg_partial_sum(reg_psum_54_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_41( .activation_in(reg_activation_54_40), .weight_in(reg_weight_53_41), .partial_sum_in(reg_psum_53_41), .reg_activation(reg_activation_54_41), .reg_weight(reg_weight_54_41), .reg_partial_sum(reg_psum_54_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_42( .activation_in(reg_activation_54_41), .weight_in(reg_weight_53_42), .partial_sum_in(reg_psum_53_42), .reg_activation(reg_activation_54_42), .reg_weight(reg_weight_54_42), .reg_partial_sum(reg_psum_54_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_43( .activation_in(reg_activation_54_42), .weight_in(reg_weight_53_43), .partial_sum_in(reg_psum_53_43), .reg_activation(reg_activation_54_43), .reg_weight(reg_weight_54_43), .reg_partial_sum(reg_psum_54_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_44( .activation_in(reg_activation_54_43), .weight_in(reg_weight_53_44), .partial_sum_in(reg_psum_53_44), .reg_activation(reg_activation_54_44), .reg_weight(reg_weight_54_44), .reg_partial_sum(reg_psum_54_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_45( .activation_in(reg_activation_54_44), .weight_in(reg_weight_53_45), .partial_sum_in(reg_psum_53_45), .reg_activation(reg_activation_54_45), .reg_weight(reg_weight_54_45), .reg_partial_sum(reg_psum_54_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_46( .activation_in(reg_activation_54_45), .weight_in(reg_weight_53_46), .partial_sum_in(reg_psum_53_46), .reg_activation(reg_activation_54_46), .reg_weight(reg_weight_54_46), .reg_partial_sum(reg_psum_54_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_47( .activation_in(reg_activation_54_46), .weight_in(reg_weight_53_47), .partial_sum_in(reg_psum_53_47), .reg_activation(reg_activation_54_47), .reg_weight(reg_weight_54_47), .reg_partial_sum(reg_psum_54_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_48( .activation_in(reg_activation_54_47), .weight_in(reg_weight_53_48), .partial_sum_in(reg_psum_53_48), .reg_activation(reg_activation_54_48), .reg_weight(reg_weight_54_48), .reg_partial_sum(reg_psum_54_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_49( .activation_in(reg_activation_54_48), .weight_in(reg_weight_53_49), .partial_sum_in(reg_psum_53_49), .reg_activation(reg_activation_54_49), .reg_weight(reg_weight_54_49), .reg_partial_sum(reg_psum_54_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_50( .activation_in(reg_activation_54_49), .weight_in(reg_weight_53_50), .partial_sum_in(reg_psum_53_50), .reg_activation(reg_activation_54_50), .reg_weight(reg_weight_54_50), .reg_partial_sum(reg_psum_54_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_51( .activation_in(reg_activation_54_50), .weight_in(reg_weight_53_51), .partial_sum_in(reg_psum_53_51), .reg_activation(reg_activation_54_51), .reg_weight(reg_weight_54_51), .reg_partial_sum(reg_psum_54_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_52( .activation_in(reg_activation_54_51), .weight_in(reg_weight_53_52), .partial_sum_in(reg_psum_53_52), .reg_activation(reg_activation_54_52), .reg_weight(reg_weight_54_52), .reg_partial_sum(reg_psum_54_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_53( .activation_in(reg_activation_54_52), .weight_in(reg_weight_53_53), .partial_sum_in(reg_psum_53_53), .reg_activation(reg_activation_54_53), .reg_weight(reg_weight_54_53), .reg_partial_sum(reg_psum_54_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_54( .activation_in(reg_activation_54_53), .weight_in(reg_weight_53_54), .partial_sum_in(reg_psum_53_54), .reg_activation(reg_activation_54_54), .reg_weight(reg_weight_54_54), .reg_partial_sum(reg_psum_54_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_55( .activation_in(reg_activation_54_54), .weight_in(reg_weight_53_55), .partial_sum_in(reg_psum_53_55), .reg_activation(reg_activation_54_55), .reg_weight(reg_weight_54_55), .reg_partial_sum(reg_psum_54_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_56( .activation_in(reg_activation_54_55), .weight_in(reg_weight_53_56), .partial_sum_in(reg_psum_53_56), .reg_activation(reg_activation_54_56), .reg_weight(reg_weight_54_56), .reg_partial_sum(reg_psum_54_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_57( .activation_in(reg_activation_54_56), .weight_in(reg_weight_53_57), .partial_sum_in(reg_psum_53_57), .reg_activation(reg_activation_54_57), .reg_weight(reg_weight_54_57), .reg_partial_sum(reg_psum_54_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_58( .activation_in(reg_activation_54_57), .weight_in(reg_weight_53_58), .partial_sum_in(reg_psum_53_58), .reg_activation(reg_activation_54_58), .reg_weight(reg_weight_54_58), .reg_partial_sum(reg_psum_54_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_59( .activation_in(reg_activation_54_58), .weight_in(reg_weight_53_59), .partial_sum_in(reg_psum_53_59), .reg_activation(reg_activation_54_59), .reg_weight(reg_weight_54_59), .reg_partial_sum(reg_psum_54_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_60( .activation_in(reg_activation_54_59), .weight_in(reg_weight_53_60), .partial_sum_in(reg_psum_53_60), .reg_activation(reg_activation_54_60), .reg_weight(reg_weight_54_60), .reg_partial_sum(reg_psum_54_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_61( .activation_in(reg_activation_54_60), .weight_in(reg_weight_53_61), .partial_sum_in(reg_psum_53_61), .reg_activation(reg_activation_54_61), .reg_weight(reg_weight_54_61), .reg_partial_sum(reg_psum_54_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_62( .activation_in(reg_activation_54_61), .weight_in(reg_weight_53_62), .partial_sum_in(reg_psum_53_62), .reg_activation(reg_activation_54_62), .reg_weight(reg_weight_54_62), .reg_partial_sum(reg_psum_54_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U54_63( .activation_in(reg_activation_54_62), .weight_in(reg_weight_53_63), .partial_sum_in(reg_psum_53_63), .reg_weight(reg_weight_54_63), .reg_partial_sum(reg_psum_54_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_0( .activation_in(in_activation_55), .weight_in(reg_weight_54_0), .partial_sum_in(reg_psum_54_0), .reg_activation(reg_activation_55_0), .reg_weight(reg_weight_55_0), .reg_partial_sum(reg_psum_55_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_1( .activation_in(reg_activation_55_0), .weight_in(reg_weight_54_1), .partial_sum_in(reg_psum_54_1), .reg_activation(reg_activation_55_1), .reg_weight(reg_weight_55_1), .reg_partial_sum(reg_psum_55_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_2( .activation_in(reg_activation_55_1), .weight_in(reg_weight_54_2), .partial_sum_in(reg_psum_54_2), .reg_activation(reg_activation_55_2), .reg_weight(reg_weight_55_2), .reg_partial_sum(reg_psum_55_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_3( .activation_in(reg_activation_55_2), .weight_in(reg_weight_54_3), .partial_sum_in(reg_psum_54_3), .reg_activation(reg_activation_55_3), .reg_weight(reg_weight_55_3), .reg_partial_sum(reg_psum_55_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_4( .activation_in(reg_activation_55_3), .weight_in(reg_weight_54_4), .partial_sum_in(reg_psum_54_4), .reg_activation(reg_activation_55_4), .reg_weight(reg_weight_55_4), .reg_partial_sum(reg_psum_55_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_5( .activation_in(reg_activation_55_4), .weight_in(reg_weight_54_5), .partial_sum_in(reg_psum_54_5), .reg_activation(reg_activation_55_5), .reg_weight(reg_weight_55_5), .reg_partial_sum(reg_psum_55_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_6( .activation_in(reg_activation_55_5), .weight_in(reg_weight_54_6), .partial_sum_in(reg_psum_54_6), .reg_activation(reg_activation_55_6), .reg_weight(reg_weight_55_6), .reg_partial_sum(reg_psum_55_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_7( .activation_in(reg_activation_55_6), .weight_in(reg_weight_54_7), .partial_sum_in(reg_psum_54_7), .reg_activation(reg_activation_55_7), .reg_weight(reg_weight_55_7), .reg_partial_sum(reg_psum_55_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_8( .activation_in(reg_activation_55_7), .weight_in(reg_weight_54_8), .partial_sum_in(reg_psum_54_8), .reg_activation(reg_activation_55_8), .reg_weight(reg_weight_55_8), .reg_partial_sum(reg_psum_55_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_9( .activation_in(reg_activation_55_8), .weight_in(reg_weight_54_9), .partial_sum_in(reg_psum_54_9), .reg_activation(reg_activation_55_9), .reg_weight(reg_weight_55_9), .reg_partial_sum(reg_psum_55_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_10( .activation_in(reg_activation_55_9), .weight_in(reg_weight_54_10), .partial_sum_in(reg_psum_54_10), .reg_activation(reg_activation_55_10), .reg_weight(reg_weight_55_10), .reg_partial_sum(reg_psum_55_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_11( .activation_in(reg_activation_55_10), .weight_in(reg_weight_54_11), .partial_sum_in(reg_psum_54_11), .reg_activation(reg_activation_55_11), .reg_weight(reg_weight_55_11), .reg_partial_sum(reg_psum_55_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_12( .activation_in(reg_activation_55_11), .weight_in(reg_weight_54_12), .partial_sum_in(reg_psum_54_12), .reg_activation(reg_activation_55_12), .reg_weight(reg_weight_55_12), .reg_partial_sum(reg_psum_55_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_13( .activation_in(reg_activation_55_12), .weight_in(reg_weight_54_13), .partial_sum_in(reg_psum_54_13), .reg_activation(reg_activation_55_13), .reg_weight(reg_weight_55_13), .reg_partial_sum(reg_psum_55_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_14( .activation_in(reg_activation_55_13), .weight_in(reg_weight_54_14), .partial_sum_in(reg_psum_54_14), .reg_activation(reg_activation_55_14), .reg_weight(reg_weight_55_14), .reg_partial_sum(reg_psum_55_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_15( .activation_in(reg_activation_55_14), .weight_in(reg_weight_54_15), .partial_sum_in(reg_psum_54_15), .reg_activation(reg_activation_55_15), .reg_weight(reg_weight_55_15), .reg_partial_sum(reg_psum_55_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_16( .activation_in(reg_activation_55_15), .weight_in(reg_weight_54_16), .partial_sum_in(reg_psum_54_16), .reg_activation(reg_activation_55_16), .reg_weight(reg_weight_55_16), .reg_partial_sum(reg_psum_55_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_17( .activation_in(reg_activation_55_16), .weight_in(reg_weight_54_17), .partial_sum_in(reg_psum_54_17), .reg_activation(reg_activation_55_17), .reg_weight(reg_weight_55_17), .reg_partial_sum(reg_psum_55_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_18( .activation_in(reg_activation_55_17), .weight_in(reg_weight_54_18), .partial_sum_in(reg_psum_54_18), .reg_activation(reg_activation_55_18), .reg_weight(reg_weight_55_18), .reg_partial_sum(reg_psum_55_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_19( .activation_in(reg_activation_55_18), .weight_in(reg_weight_54_19), .partial_sum_in(reg_psum_54_19), .reg_activation(reg_activation_55_19), .reg_weight(reg_weight_55_19), .reg_partial_sum(reg_psum_55_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_20( .activation_in(reg_activation_55_19), .weight_in(reg_weight_54_20), .partial_sum_in(reg_psum_54_20), .reg_activation(reg_activation_55_20), .reg_weight(reg_weight_55_20), .reg_partial_sum(reg_psum_55_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_21( .activation_in(reg_activation_55_20), .weight_in(reg_weight_54_21), .partial_sum_in(reg_psum_54_21), .reg_activation(reg_activation_55_21), .reg_weight(reg_weight_55_21), .reg_partial_sum(reg_psum_55_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_22( .activation_in(reg_activation_55_21), .weight_in(reg_weight_54_22), .partial_sum_in(reg_psum_54_22), .reg_activation(reg_activation_55_22), .reg_weight(reg_weight_55_22), .reg_partial_sum(reg_psum_55_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_23( .activation_in(reg_activation_55_22), .weight_in(reg_weight_54_23), .partial_sum_in(reg_psum_54_23), .reg_activation(reg_activation_55_23), .reg_weight(reg_weight_55_23), .reg_partial_sum(reg_psum_55_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_24( .activation_in(reg_activation_55_23), .weight_in(reg_weight_54_24), .partial_sum_in(reg_psum_54_24), .reg_activation(reg_activation_55_24), .reg_weight(reg_weight_55_24), .reg_partial_sum(reg_psum_55_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_25( .activation_in(reg_activation_55_24), .weight_in(reg_weight_54_25), .partial_sum_in(reg_psum_54_25), .reg_activation(reg_activation_55_25), .reg_weight(reg_weight_55_25), .reg_partial_sum(reg_psum_55_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_26( .activation_in(reg_activation_55_25), .weight_in(reg_weight_54_26), .partial_sum_in(reg_psum_54_26), .reg_activation(reg_activation_55_26), .reg_weight(reg_weight_55_26), .reg_partial_sum(reg_psum_55_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_27( .activation_in(reg_activation_55_26), .weight_in(reg_weight_54_27), .partial_sum_in(reg_psum_54_27), .reg_activation(reg_activation_55_27), .reg_weight(reg_weight_55_27), .reg_partial_sum(reg_psum_55_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_28( .activation_in(reg_activation_55_27), .weight_in(reg_weight_54_28), .partial_sum_in(reg_psum_54_28), .reg_activation(reg_activation_55_28), .reg_weight(reg_weight_55_28), .reg_partial_sum(reg_psum_55_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_29( .activation_in(reg_activation_55_28), .weight_in(reg_weight_54_29), .partial_sum_in(reg_psum_54_29), .reg_activation(reg_activation_55_29), .reg_weight(reg_weight_55_29), .reg_partial_sum(reg_psum_55_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_30( .activation_in(reg_activation_55_29), .weight_in(reg_weight_54_30), .partial_sum_in(reg_psum_54_30), .reg_activation(reg_activation_55_30), .reg_weight(reg_weight_55_30), .reg_partial_sum(reg_psum_55_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_31( .activation_in(reg_activation_55_30), .weight_in(reg_weight_54_31), .partial_sum_in(reg_psum_54_31), .reg_activation(reg_activation_55_31), .reg_weight(reg_weight_55_31), .reg_partial_sum(reg_psum_55_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_32( .activation_in(reg_activation_55_31), .weight_in(reg_weight_54_32), .partial_sum_in(reg_psum_54_32), .reg_activation(reg_activation_55_32), .reg_weight(reg_weight_55_32), .reg_partial_sum(reg_psum_55_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_33( .activation_in(reg_activation_55_32), .weight_in(reg_weight_54_33), .partial_sum_in(reg_psum_54_33), .reg_activation(reg_activation_55_33), .reg_weight(reg_weight_55_33), .reg_partial_sum(reg_psum_55_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_34( .activation_in(reg_activation_55_33), .weight_in(reg_weight_54_34), .partial_sum_in(reg_psum_54_34), .reg_activation(reg_activation_55_34), .reg_weight(reg_weight_55_34), .reg_partial_sum(reg_psum_55_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_35( .activation_in(reg_activation_55_34), .weight_in(reg_weight_54_35), .partial_sum_in(reg_psum_54_35), .reg_activation(reg_activation_55_35), .reg_weight(reg_weight_55_35), .reg_partial_sum(reg_psum_55_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_36( .activation_in(reg_activation_55_35), .weight_in(reg_weight_54_36), .partial_sum_in(reg_psum_54_36), .reg_activation(reg_activation_55_36), .reg_weight(reg_weight_55_36), .reg_partial_sum(reg_psum_55_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_37( .activation_in(reg_activation_55_36), .weight_in(reg_weight_54_37), .partial_sum_in(reg_psum_54_37), .reg_activation(reg_activation_55_37), .reg_weight(reg_weight_55_37), .reg_partial_sum(reg_psum_55_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_38( .activation_in(reg_activation_55_37), .weight_in(reg_weight_54_38), .partial_sum_in(reg_psum_54_38), .reg_activation(reg_activation_55_38), .reg_weight(reg_weight_55_38), .reg_partial_sum(reg_psum_55_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_39( .activation_in(reg_activation_55_38), .weight_in(reg_weight_54_39), .partial_sum_in(reg_psum_54_39), .reg_activation(reg_activation_55_39), .reg_weight(reg_weight_55_39), .reg_partial_sum(reg_psum_55_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_40( .activation_in(reg_activation_55_39), .weight_in(reg_weight_54_40), .partial_sum_in(reg_psum_54_40), .reg_activation(reg_activation_55_40), .reg_weight(reg_weight_55_40), .reg_partial_sum(reg_psum_55_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_41( .activation_in(reg_activation_55_40), .weight_in(reg_weight_54_41), .partial_sum_in(reg_psum_54_41), .reg_activation(reg_activation_55_41), .reg_weight(reg_weight_55_41), .reg_partial_sum(reg_psum_55_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_42( .activation_in(reg_activation_55_41), .weight_in(reg_weight_54_42), .partial_sum_in(reg_psum_54_42), .reg_activation(reg_activation_55_42), .reg_weight(reg_weight_55_42), .reg_partial_sum(reg_psum_55_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_43( .activation_in(reg_activation_55_42), .weight_in(reg_weight_54_43), .partial_sum_in(reg_psum_54_43), .reg_activation(reg_activation_55_43), .reg_weight(reg_weight_55_43), .reg_partial_sum(reg_psum_55_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_44( .activation_in(reg_activation_55_43), .weight_in(reg_weight_54_44), .partial_sum_in(reg_psum_54_44), .reg_activation(reg_activation_55_44), .reg_weight(reg_weight_55_44), .reg_partial_sum(reg_psum_55_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_45( .activation_in(reg_activation_55_44), .weight_in(reg_weight_54_45), .partial_sum_in(reg_psum_54_45), .reg_activation(reg_activation_55_45), .reg_weight(reg_weight_55_45), .reg_partial_sum(reg_psum_55_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_46( .activation_in(reg_activation_55_45), .weight_in(reg_weight_54_46), .partial_sum_in(reg_psum_54_46), .reg_activation(reg_activation_55_46), .reg_weight(reg_weight_55_46), .reg_partial_sum(reg_psum_55_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_47( .activation_in(reg_activation_55_46), .weight_in(reg_weight_54_47), .partial_sum_in(reg_psum_54_47), .reg_activation(reg_activation_55_47), .reg_weight(reg_weight_55_47), .reg_partial_sum(reg_psum_55_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_48( .activation_in(reg_activation_55_47), .weight_in(reg_weight_54_48), .partial_sum_in(reg_psum_54_48), .reg_activation(reg_activation_55_48), .reg_weight(reg_weight_55_48), .reg_partial_sum(reg_psum_55_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_49( .activation_in(reg_activation_55_48), .weight_in(reg_weight_54_49), .partial_sum_in(reg_psum_54_49), .reg_activation(reg_activation_55_49), .reg_weight(reg_weight_55_49), .reg_partial_sum(reg_psum_55_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_50( .activation_in(reg_activation_55_49), .weight_in(reg_weight_54_50), .partial_sum_in(reg_psum_54_50), .reg_activation(reg_activation_55_50), .reg_weight(reg_weight_55_50), .reg_partial_sum(reg_psum_55_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_51( .activation_in(reg_activation_55_50), .weight_in(reg_weight_54_51), .partial_sum_in(reg_psum_54_51), .reg_activation(reg_activation_55_51), .reg_weight(reg_weight_55_51), .reg_partial_sum(reg_psum_55_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_52( .activation_in(reg_activation_55_51), .weight_in(reg_weight_54_52), .partial_sum_in(reg_psum_54_52), .reg_activation(reg_activation_55_52), .reg_weight(reg_weight_55_52), .reg_partial_sum(reg_psum_55_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_53( .activation_in(reg_activation_55_52), .weight_in(reg_weight_54_53), .partial_sum_in(reg_psum_54_53), .reg_activation(reg_activation_55_53), .reg_weight(reg_weight_55_53), .reg_partial_sum(reg_psum_55_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_54( .activation_in(reg_activation_55_53), .weight_in(reg_weight_54_54), .partial_sum_in(reg_psum_54_54), .reg_activation(reg_activation_55_54), .reg_weight(reg_weight_55_54), .reg_partial_sum(reg_psum_55_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_55( .activation_in(reg_activation_55_54), .weight_in(reg_weight_54_55), .partial_sum_in(reg_psum_54_55), .reg_activation(reg_activation_55_55), .reg_weight(reg_weight_55_55), .reg_partial_sum(reg_psum_55_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_56( .activation_in(reg_activation_55_55), .weight_in(reg_weight_54_56), .partial_sum_in(reg_psum_54_56), .reg_activation(reg_activation_55_56), .reg_weight(reg_weight_55_56), .reg_partial_sum(reg_psum_55_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_57( .activation_in(reg_activation_55_56), .weight_in(reg_weight_54_57), .partial_sum_in(reg_psum_54_57), .reg_activation(reg_activation_55_57), .reg_weight(reg_weight_55_57), .reg_partial_sum(reg_psum_55_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_58( .activation_in(reg_activation_55_57), .weight_in(reg_weight_54_58), .partial_sum_in(reg_psum_54_58), .reg_activation(reg_activation_55_58), .reg_weight(reg_weight_55_58), .reg_partial_sum(reg_psum_55_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_59( .activation_in(reg_activation_55_58), .weight_in(reg_weight_54_59), .partial_sum_in(reg_psum_54_59), .reg_activation(reg_activation_55_59), .reg_weight(reg_weight_55_59), .reg_partial_sum(reg_psum_55_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_60( .activation_in(reg_activation_55_59), .weight_in(reg_weight_54_60), .partial_sum_in(reg_psum_54_60), .reg_activation(reg_activation_55_60), .reg_weight(reg_weight_55_60), .reg_partial_sum(reg_psum_55_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_61( .activation_in(reg_activation_55_60), .weight_in(reg_weight_54_61), .partial_sum_in(reg_psum_54_61), .reg_activation(reg_activation_55_61), .reg_weight(reg_weight_55_61), .reg_partial_sum(reg_psum_55_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_62( .activation_in(reg_activation_55_61), .weight_in(reg_weight_54_62), .partial_sum_in(reg_psum_54_62), .reg_activation(reg_activation_55_62), .reg_weight(reg_weight_55_62), .reg_partial_sum(reg_psum_55_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U55_63( .activation_in(reg_activation_55_62), .weight_in(reg_weight_54_63), .partial_sum_in(reg_psum_54_63), .reg_weight(reg_weight_55_63), .reg_partial_sum(reg_psum_55_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_0( .activation_in(in_activation_56), .weight_in(reg_weight_55_0), .partial_sum_in(reg_psum_55_0), .reg_activation(reg_activation_56_0), .reg_weight(reg_weight_56_0), .reg_partial_sum(reg_psum_56_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_1( .activation_in(reg_activation_56_0), .weight_in(reg_weight_55_1), .partial_sum_in(reg_psum_55_1), .reg_activation(reg_activation_56_1), .reg_weight(reg_weight_56_1), .reg_partial_sum(reg_psum_56_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_2( .activation_in(reg_activation_56_1), .weight_in(reg_weight_55_2), .partial_sum_in(reg_psum_55_2), .reg_activation(reg_activation_56_2), .reg_weight(reg_weight_56_2), .reg_partial_sum(reg_psum_56_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_3( .activation_in(reg_activation_56_2), .weight_in(reg_weight_55_3), .partial_sum_in(reg_psum_55_3), .reg_activation(reg_activation_56_3), .reg_weight(reg_weight_56_3), .reg_partial_sum(reg_psum_56_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_4( .activation_in(reg_activation_56_3), .weight_in(reg_weight_55_4), .partial_sum_in(reg_psum_55_4), .reg_activation(reg_activation_56_4), .reg_weight(reg_weight_56_4), .reg_partial_sum(reg_psum_56_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_5( .activation_in(reg_activation_56_4), .weight_in(reg_weight_55_5), .partial_sum_in(reg_psum_55_5), .reg_activation(reg_activation_56_5), .reg_weight(reg_weight_56_5), .reg_partial_sum(reg_psum_56_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_6( .activation_in(reg_activation_56_5), .weight_in(reg_weight_55_6), .partial_sum_in(reg_psum_55_6), .reg_activation(reg_activation_56_6), .reg_weight(reg_weight_56_6), .reg_partial_sum(reg_psum_56_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_7( .activation_in(reg_activation_56_6), .weight_in(reg_weight_55_7), .partial_sum_in(reg_psum_55_7), .reg_activation(reg_activation_56_7), .reg_weight(reg_weight_56_7), .reg_partial_sum(reg_psum_56_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_8( .activation_in(reg_activation_56_7), .weight_in(reg_weight_55_8), .partial_sum_in(reg_psum_55_8), .reg_activation(reg_activation_56_8), .reg_weight(reg_weight_56_8), .reg_partial_sum(reg_psum_56_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_9( .activation_in(reg_activation_56_8), .weight_in(reg_weight_55_9), .partial_sum_in(reg_psum_55_9), .reg_activation(reg_activation_56_9), .reg_weight(reg_weight_56_9), .reg_partial_sum(reg_psum_56_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_10( .activation_in(reg_activation_56_9), .weight_in(reg_weight_55_10), .partial_sum_in(reg_psum_55_10), .reg_activation(reg_activation_56_10), .reg_weight(reg_weight_56_10), .reg_partial_sum(reg_psum_56_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_11( .activation_in(reg_activation_56_10), .weight_in(reg_weight_55_11), .partial_sum_in(reg_psum_55_11), .reg_activation(reg_activation_56_11), .reg_weight(reg_weight_56_11), .reg_partial_sum(reg_psum_56_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_12( .activation_in(reg_activation_56_11), .weight_in(reg_weight_55_12), .partial_sum_in(reg_psum_55_12), .reg_activation(reg_activation_56_12), .reg_weight(reg_weight_56_12), .reg_partial_sum(reg_psum_56_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_13( .activation_in(reg_activation_56_12), .weight_in(reg_weight_55_13), .partial_sum_in(reg_psum_55_13), .reg_activation(reg_activation_56_13), .reg_weight(reg_weight_56_13), .reg_partial_sum(reg_psum_56_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_14( .activation_in(reg_activation_56_13), .weight_in(reg_weight_55_14), .partial_sum_in(reg_psum_55_14), .reg_activation(reg_activation_56_14), .reg_weight(reg_weight_56_14), .reg_partial_sum(reg_psum_56_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_15( .activation_in(reg_activation_56_14), .weight_in(reg_weight_55_15), .partial_sum_in(reg_psum_55_15), .reg_activation(reg_activation_56_15), .reg_weight(reg_weight_56_15), .reg_partial_sum(reg_psum_56_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_16( .activation_in(reg_activation_56_15), .weight_in(reg_weight_55_16), .partial_sum_in(reg_psum_55_16), .reg_activation(reg_activation_56_16), .reg_weight(reg_weight_56_16), .reg_partial_sum(reg_psum_56_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_17( .activation_in(reg_activation_56_16), .weight_in(reg_weight_55_17), .partial_sum_in(reg_psum_55_17), .reg_activation(reg_activation_56_17), .reg_weight(reg_weight_56_17), .reg_partial_sum(reg_psum_56_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_18( .activation_in(reg_activation_56_17), .weight_in(reg_weight_55_18), .partial_sum_in(reg_psum_55_18), .reg_activation(reg_activation_56_18), .reg_weight(reg_weight_56_18), .reg_partial_sum(reg_psum_56_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_19( .activation_in(reg_activation_56_18), .weight_in(reg_weight_55_19), .partial_sum_in(reg_psum_55_19), .reg_activation(reg_activation_56_19), .reg_weight(reg_weight_56_19), .reg_partial_sum(reg_psum_56_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_20( .activation_in(reg_activation_56_19), .weight_in(reg_weight_55_20), .partial_sum_in(reg_psum_55_20), .reg_activation(reg_activation_56_20), .reg_weight(reg_weight_56_20), .reg_partial_sum(reg_psum_56_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_21( .activation_in(reg_activation_56_20), .weight_in(reg_weight_55_21), .partial_sum_in(reg_psum_55_21), .reg_activation(reg_activation_56_21), .reg_weight(reg_weight_56_21), .reg_partial_sum(reg_psum_56_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_22( .activation_in(reg_activation_56_21), .weight_in(reg_weight_55_22), .partial_sum_in(reg_psum_55_22), .reg_activation(reg_activation_56_22), .reg_weight(reg_weight_56_22), .reg_partial_sum(reg_psum_56_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_23( .activation_in(reg_activation_56_22), .weight_in(reg_weight_55_23), .partial_sum_in(reg_psum_55_23), .reg_activation(reg_activation_56_23), .reg_weight(reg_weight_56_23), .reg_partial_sum(reg_psum_56_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_24( .activation_in(reg_activation_56_23), .weight_in(reg_weight_55_24), .partial_sum_in(reg_psum_55_24), .reg_activation(reg_activation_56_24), .reg_weight(reg_weight_56_24), .reg_partial_sum(reg_psum_56_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_25( .activation_in(reg_activation_56_24), .weight_in(reg_weight_55_25), .partial_sum_in(reg_psum_55_25), .reg_activation(reg_activation_56_25), .reg_weight(reg_weight_56_25), .reg_partial_sum(reg_psum_56_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_26( .activation_in(reg_activation_56_25), .weight_in(reg_weight_55_26), .partial_sum_in(reg_psum_55_26), .reg_activation(reg_activation_56_26), .reg_weight(reg_weight_56_26), .reg_partial_sum(reg_psum_56_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_27( .activation_in(reg_activation_56_26), .weight_in(reg_weight_55_27), .partial_sum_in(reg_psum_55_27), .reg_activation(reg_activation_56_27), .reg_weight(reg_weight_56_27), .reg_partial_sum(reg_psum_56_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_28( .activation_in(reg_activation_56_27), .weight_in(reg_weight_55_28), .partial_sum_in(reg_psum_55_28), .reg_activation(reg_activation_56_28), .reg_weight(reg_weight_56_28), .reg_partial_sum(reg_psum_56_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_29( .activation_in(reg_activation_56_28), .weight_in(reg_weight_55_29), .partial_sum_in(reg_psum_55_29), .reg_activation(reg_activation_56_29), .reg_weight(reg_weight_56_29), .reg_partial_sum(reg_psum_56_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_30( .activation_in(reg_activation_56_29), .weight_in(reg_weight_55_30), .partial_sum_in(reg_psum_55_30), .reg_activation(reg_activation_56_30), .reg_weight(reg_weight_56_30), .reg_partial_sum(reg_psum_56_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_31( .activation_in(reg_activation_56_30), .weight_in(reg_weight_55_31), .partial_sum_in(reg_psum_55_31), .reg_activation(reg_activation_56_31), .reg_weight(reg_weight_56_31), .reg_partial_sum(reg_psum_56_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_32( .activation_in(reg_activation_56_31), .weight_in(reg_weight_55_32), .partial_sum_in(reg_psum_55_32), .reg_activation(reg_activation_56_32), .reg_weight(reg_weight_56_32), .reg_partial_sum(reg_psum_56_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_33( .activation_in(reg_activation_56_32), .weight_in(reg_weight_55_33), .partial_sum_in(reg_psum_55_33), .reg_activation(reg_activation_56_33), .reg_weight(reg_weight_56_33), .reg_partial_sum(reg_psum_56_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_34( .activation_in(reg_activation_56_33), .weight_in(reg_weight_55_34), .partial_sum_in(reg_psum_55_34), .reg_activation(reg_activation_56_34), .reg_weight(reg_weight_56_34), .reg_partial_sum(reg_psum_56_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_35( .activation_in(reg_activation_56_34), .weight_in(reg_weight_55_35), .partial_sum_in(reg_psum_55_35), .reg_activation(reg_activation_56_35), .reg_weight(reg_weight_56_35), .reg_partial_sum(reg_psum_56_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_36( .activation_in(reg_activation_56_35), .weight_in(reg_weight_55_36), .partial_sum_in(reg_psum_55_36), .reg_activation(reg_activation_56_36), .reg_weight(reg_weight_56_36), .reg_partial_sum(reg_psum_56_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_37( .activation_in(reg_activation_56_36), .weight_in(reg_weight_55_37), .partial_sum_in(reg_psum_55_37), .reg_activation(reg_activation_56_37), .reg_weight(reg_weight_56_37), .reg_partial_sum(reg_psum_56_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_38( .activation_in(reg_activation_56_37), .weight_in(reg_weight_55_38), .partial_sum_in(reg_psum_55_38), .reg_activation(reg_activation_56_38), .reg_weight(reg_weight_56_38), .reg_partial_sum(reg_psum_56_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_39( .activation_in(reg_activation_56_38), .weight_in(reg_weight_55_39), .partial_sum_in(reg_psum_55_39), .reg_activation(reg_activation_56_39), .reg_weight(reg_weight_56_39), .reg_partial_sum(reg_psum_56_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_40( .activation_in(reg_activation_56_39), .weight_in(reg_weight_55_40), .partial_sum_in(reg_psum_55_40), .reg_activation(reg_activation_56_40), .reg_weight(reg_weight_56_40), .reg_partial_sum(reg_psum_56_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_41( .activation_in(reg_activation_56_40), .weight_in(reg_weight_55_41), .partial_sum_in(reg_psum_55_41), .reg_activation(reg_activation_56_41), .reg_weight(reg_weight_56_41), .reg_partial_sum(reg_psum_56_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_42( .activation_in(reg_activation_56_41), .weight_in(reg_weight_55_42), .partial_sum_in(reg_psum_55_42), .reg_activation(reg_activation_56_42), .reg_weight(reg_weight_56_42), .reg_partial_sum(reg_psum_56_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_43( .activation_in(reg_activation_56_42), .weight_in(reg_weight_55_43), .partial_sum_in(reg_psum_55_43), .reg_activation(reg_activation_56_43), .reg_weight(reg_weight_56_43), .reg_partial_sum(reg_psum_56_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_44( .activation_in(reg_activation_56_43), .weight_in(reg_weight_55_44), .partial_sum_in(reg_psum_55_44), .reg_activation(reg_activation_56_44), .reg_weight(reg_weight_56_44), .reg_partial_sum(reg_psum_56_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_45( .activation_in(reg_activation_56_44), .weight_in(reg_weight_55_45), .partial_sum_in(reg_psum_55_45), .reg_activation(reg_activation_56_45), .reg_weight(reg_weight_56_45), .reg_partial_sum(reg_psum_56_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_46( .activation_in(reg_activation_56_45), .weight_in(reg_weight_55_46), .partial_sum_in(reg_psum_55_46), .reg_activation(reg_activation_56_46), .reg_weight(reg_weight_56_46), .reg_partial_sum(reg_psum_56_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_47( .activation_in(reg_activation_56_46), .weight_in(reg_weight_55_47), .partial_sum_in(reg_psum_55_47), .reg_activation(reg_activation_56_47), .reg_weight(reg_weight_56_47), .reg_partial_sum(reg_psum_56_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_48( .activation_in(reg_activation_56_47), .weight_in(reg_weight_55_48), .partial_sum_in(reg_psum_55_48), .reg_activation(reg_activation_56_48), .reg_weight(reg_weight_56_48), .reg_partial_sum(reg_psum_56_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_49( .activation_in(reg_activation_56_48), .weight_in(reg_weight_55_49), .partial_sum_in(reg_psum_55_49), .reg_activation(reg_activation_56_49), .reg_weight(reg_weight_56_49), .reg_partial_sum(reg_psum_56_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_50( .activation_in(reg_activation_56_49), .weight_in(reg_weight_55_50), .partial_sum_in(reg_psum_55_50), .reg_activation(reg_activation_56_50), .reg_weight(reg_weight_56_50), .reg_partial_sum(reg_psum_56_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_51( .activation_in(reg_activation_56_50), .weight_in(reg_weight_55_51), .partial_sum_in(reg_psum_55_51), .reg_activation(reg_activation_56_51), .reg_weight(reg_weight_56_51), .reg_partial_sum(reg_psum_56_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_52( .activation_in(reg_activation_56_51), .weight_in(reg_weight_55_52), .partial_sum_in(reg_psum_55_52), .reg_activation(reg_activation_56_52), .reg_weight(reg_weight_56_52), .reg_partial_sum(reg_psum_56_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_53( .activation_in(reg_activation_56_52), .weight_in(reg_weight_55_53), .partial_sum_in(reg_psum_55_53), .reg_activation(reg_activation_56_53), .reg_weight(reg_weight_56_53), .reg_partial_sum(reg_psum_56_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_54( .activation_in(reg_activation_56_53), .weight_in(reg_weight_55_54), .partial_sum_in(reg_psum_55_54), .reg_activation(reg_activation_56_54), .reg_weight(reg_weight_56_54), .reg_partial_sum(reg_psum_56_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_55( .activation_in(reg_activation_56_54), .weight_in(reg_weight_55_55), .partial_sum_in(reg_psum_55_55), .reg_activation(reg_activation_56_55), .reg_weight(reg_weight_56_55), .reg_partial_sum(reg_psum_56_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_56( .activation_in(reg_activation_56_55), .weight_in(reg_weight_55_56), .partial_sum_in(reg_psum_55_56), .reg_activation(reg_activation_56_56), .reg_weight(reg_weight_56_56), .reg_partial_sum(reg_psum_56_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_57( .activation_in(reg_activation_56_56), .weight_in(reg_weight_55_57), .partial_sum_in(reg_psum_55_57), .reg_activation(reg_activation_56_57), .reg_weight(reg_weight_56_57), .reg_partial_sum(reg_psum_56_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_58( .activation_in(reg_activation_56_57), .weight_in(reg_weight_55_58), .partial_sum_in(reg_psum_55_58), .reg_activation(reg_activation_56_58), .reg_weight(reg_weight_56_58), .reg_partial_sum(reg_psum_56_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_59( .activation_in(reg_activation_56_58), .weight_in(reg_weight_55_59), .partial_sum_in(reg_psum_55_59), .reg_activation(reg_activation_56_59), .reg_weight(reg_weight_56_59), .reg_partial_sum(reg_psum_56_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_60( .activation_in(reg_activation_56_59), .weight_in(reg_weight_55_60), .partial_sum_in(reg_psum_55_60), .reg_activation(reg_activation_56_60), .reg_weight(reg_weight_56_60), .reg_partial_sum(reg_psum_56_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_61( .activation_in(reg_activation_56_60), .weight_in(reg_weight_55_61), .partial_sum_in(reg_psum_55_61), .reg_activation(reg_activation_56_61), .reg_weight(reg_weight_56_61), .reg_partial_sum(reg_psum_56_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_62( .activation_in(reg_activation_56_61), .weight_in(reg_weight_55_62), .partial_sum_in(reg_psum_55_62), .reg_activation(reg_activation_56_62), .reg_weight(reg_weight_56_62), .reg_partial_sum(reg_psum_56_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U56_63( .activation_in(reg_activation_56_62), .weight_in(reg_weight_55_63), .partial_sum_in(reg_psum_55_63), .reg_weight(reg_weight_56_63), .reg_partial_sum(reg_psum_56_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_0( .activation_in(in_activation_57), .weight_in(reg_weight_56_0), .partial_sum_in(reg_psum_56_0), .reg_activation(reg_activation_57_0), .reg_weight(reg_weight_57_0), .reg_partial_sum(reg_psum_57_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_1( .activation_in(reg_activation_57_0), .weight_in(reg_weight_56_1), .partial_sum_in(reg_psum_56_1), .reg_activation(reg_activation_57_1), .reg_weight(reg_weight_57_1), .reg_partial_sum(reg_psum_57_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_2( .activation_in(reg_activation_57_1), .weight_in(reg_weight_56_2), .partial_sum_in(reg_psum_56_2), .reg_activation(reg_activation_57_2), .reg_weight(reg_weight_57_2), .reg_partial_sum(reg_psum_57_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_3( .activation_in(reg_activation_57_2), .weight_in(reg_weight_56_3), .partial_sum_in(reg_psum_56_3), .reg_activation(reg_activation_57_3), .reg_weight(reg_weight_57_3), .reg_partial_sum(reg_psum_57_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_4( .activation_in(reg_activation_57_3), .weight_in(reg_weight_56_4), .partial_sum_in(reg_psum_56_4), .reg_activation(reg_activation_57_4), .reg_weight(reg_weight_57_4), .reg_partial_sum(reg_psum_57_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_5( .activation_in(reg_activation_57_4), .weight_in(reg_weight_56_5), .partial_sum_in(reg_psum_56_5), .reg_activation(reg_activation_57_5), .reg_weight(reg_weight_57_5), .reg_partial_sum(reg_psum_57_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_6( .activation_in(reg_activation_57_5), .weight_in(reg_weight_56_6), .partial_sum_in(reg_psum_56_6), .reg_activation(reg_activation_57_6), .reg_weight(reg_weight_57_6), .reg_partial_sum(reg_psum_57_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_7( .activation_in(reg_activation_57_6), .weight_in(reg_weight_56_7), .partial_sum_in(reg_psum_56_7), .reg_activation(reg_activation_57_7), .reg_weight(reg_weight_57_7), .reg_partial_sum(reg_psum_57_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_8( .activation_in(reg_activation_57_7), .weight_in(reg_weight_56_8), .partial_sum_in(reg_psum_56_8), .reg_activation(reg_activation_57_8), .reg_weight(reg_weight_57_8), .reg_partial_sum(reg_psum_57_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_9( .activation_in(reg_activation_57_8), .weight_in(reg_weight_56_9), .partial_sum_in(reg_psum_56_9), .reg_activation(reg_activation_57_9), .reg_weight(reg_weight_57_9), .reg_partial_sum(reg_psum_57_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_10( .activation_in(reg_activation_57_9), .weight_in(reg_weight_56_10), .partial_sum_in(reg_psum_56_10), .reg_activation(reg_activation_57_10), .reg_weight(reg_weight_57_10), .reg_partial_sum(reg_psum_57_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_11( .activation_in(reg_activation_57_10), .weight_in(reg_weight_56_11), .partial_sum_in(reg_psum_56_11), .reg_activation(reg_activation_57_11), .reg_weight(reg_weight_57_11), .reg_partial_sum(reg_psum_57_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_12( .activation_in(reg_activation_57_11), .weight_in(reg_weight_56_12), .partial_sum_in(reg_psum_56_12), .reg_activation(reg_activation_57_12), .reg_weight(reg_weight_57_12), .reg_partial_sum(reg_psum_57_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_13( .activation_in(reg_activation_57_12), .weight_in(reg_weight_56_13), .partial_sum_in(reg_psum_56_13), .reg_activation(reg_activation_57_13), .reg_weight(reg_weight_57_13), .reg_partial_sum(reg_psum_57_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_14( .activation_in(reg_activation_57_13), .weight_in(reg_weight_56_14), .partial_sum_in(reg_psum_56_14), .reg_activation(reg_activation_57_14), .reg_weight(reg_weight_57_14), .reg_partial_sum(reg_psum_57_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_15( .activation_in(reg_activation_57_14), .weight_in(reg_weight_56_15), .partial_sum_in(reg_psum_56_15), .reg_activation(reg_activation_57_15), .reg_weight(reg_weight_57_15), .reg_partial_sum(reg_psum_57_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_16( .activation_in(reg_activation_57_15), .weight_in(reg_weight_56_16), .partial_sum_in(reg_psum_56_16), .reg_activation(reg_activation_57_16), .reg_weight(reg_weight_57_16), .reg_partial_sum(reg_psum_57_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_17( .activation_in(reg_activation_57_16), .weight_in(reg_weight_56_17), .partial_sum_in(reg_psum_56_17), .reg_activation(reg_activation_57_17), .reg_weight(reg_weight_57_17), .reg_partial_sum(reg_psum_57_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_18( .activation_in(reg_activation_57_17), .weight_in(reg_weight_56_18), .partial_sum_in(reg_psum_56_18), .reg_activation(reg_activation_57_18), .reg_weight(reg_weight_57_18), .reg_partial_sum(reg_psum_57_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_19( .activation_in(reg_activation_57_18), .weight_in(reg_weight_56_19), .partial_sum_in(reg_psum_56_19), .reg_activation(reg_activation_57_19), .reg_weight(reg_weight_57_19), .reg_partial_sum(reg_psum_57_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_20( .activation_in(reg_activation_57_19), .weight_in(reg_weight_56_20), .partial_sum_in(reg_psum_56_20), .reg_activation(reg_activation_57_20), .reg_weight(reg_weight_57_20), .reg_partial_sum(reg_psum_57_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_21( .activation_in(reg_activation_57_20), .weight_in(reg_weight_56_21), .partial_sum_in(reg_psum_56_21), .reg_activation(reg_activation_57_21), .reg_weight(reg_weight_57_21), .reg_partial_sum(reg_psum_57_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_22( .activation_in(reg_activation_57_21), .weight_in(reg_weight_56_22), .partial_sum_in(reg_psum_56_22), .reg_activation(reg_activation_57_22), .reg_weight(reg_weight_57_22), .reg_partial_sum(reg_psum_57_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_23( .activation_in(reg_activation_57_22), .weight_in(reg_weight_56_23), .partial_sum_in(reg_psum_56_23), .reg_activation(reg_activation_57_23), .reg_weight(reg_weight_57_23), .reg_partial_sum(reg_psum_57_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_24( .activation_in(reg_activation_57_23), .weight_in(reg_weight_56_24), .partial_sum_in(reg_psum_56_24), .reg_activation(reg_activation_57_24), .reg_weight(reg_weight_57_24), .reg_partial_sum(reg_psum_57_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_25( .activation_in(reg_activation_57_24), .weight_in(reg_weight_56_25), .partial_sum_in(reg_psum_56_25), .reg_activation(reg_activation_57_25), .reg_weight(reg_weight_57_25), .reg_partial_sum(reg_psum_57_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_26( .activation_in(reg_activation_57_25), .weight_in(reg_weight_56_26), .partial_sum_in(reg_psum_56_26), .reg_activation(reg_activation_57_26), .reg_weight(reg_weight_57_26), .reg_partial_sum(reg_psum_57_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_27( .activation_in(reg_activation_57_26), .weight_in(reg_weight_56_27), .partial_sum_in(reg_psum_56_27), .reg_activation(reg_activation_57_27), .reg_weight(reg_weight_57_27), .reg_partial_sum(reg_psum_57_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_28( .activation_in(reg_activation_57_27), .weight_in(reg_weight_56_28), .partial_sum_in(reg_psum_56_28), .reg_activation(reg_activation_57_28), .reg_weight(reg_weight_57_28), .reg_partial_sum(reg_psum_57_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_29( .activation_in(reg_activation_57_28), .weight_in(reg_weight_56_29), .partial_sum_in(reg_psum_56_29), .reg_activation(reg_activation_57_29), .reg_weight(reg_weight_57_29), .reg_partial_sum(reg_psum_57_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_30( .activation_in(reg_activation_57_29), .weight_in(reg_weight_56_30), .partial_sum_in(reg_psum_56_30), .reg_activation(reg_activation_57_30), .reg_weight(reg_weight_57_30), .reg_partial_sum(reg_psum_57_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_31( .activation_in(reg_activation_57_30), .weight_in(reg_weight_56_31), .partial_sum_in(reg_psum_56_31), .reg_activation(reg_activation_57_31), .reg_weight(reg_weight_57_31), .reg_partial_sum(reg_psum_57_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_32( .activation_in(reg_activation_57_31), .weight_in(reg_weight_56_32), .partial_sum_in(reg_psum_56_32), .reg_activation(reg_activation_57_32), .reg_weight(reg_weight_57_32), .reg_partial_sum(reg_psum_57_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_33( .activation_in(reg_activation_57_32), .weight_in(reg_weight_56_33), .partial_sum_in(reg_psum_56_33), .reg_activation(reg_activation_57_33), .reg_weight(reg_weight_57_33), .reg_partial_sum(reg_psum_57_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_34( .activation_in(reg_activation_57_33), .weight_in(reg_weight_56_34), .partial_sum_in(reg_psum_56_34), .reg_activation(reg_activation_57_34), .reg_weight(reg_weight_57_34), .reg_partial_sum(reg_psum_57_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_35( .activation_in(reg_activation_57_34), .weight_in(reg_weight_56_35), .partial_sum_in(reg_psum_56_35), .reg_activation(reg_activation_57_35), .reg_weight(reg_weight_57_35), .reg_partial_sum(reg_psum_57_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_36( .activation_in(reg_activation_57_35), .weight_in(reg_weight_56_36), .partial_sum_in(reg_psum_56_36), .reg_activation(reg_activation_57_36), .reg_weight(reg_weight_57_36), .reg_partial_sum(reg_psum_57_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_37( .activation_in(reg_activation_57_36), .weight_in(reg_weight_56_37), .partial_sum_in(reg_psum_56_37), .reg_activation(reg_activation_57_37), .reg_weight(reg_weight_57_37), .reg_partial_sum(reg_psum_57_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_38( .activation_in(reg_activation_57_37), .weight_in(reg_weight_56_38), .partial_sum_in(reg_psum_56_38), .reg_activation(reg_activation_57_38), .reg_weight(reg_weight_57_38), .reg_partial_sum(reg_psum_57_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_39( .activation_in(reg_activation_57_38), .weight_in(reg_weight_56_39), .partial_sum_in(reg_psum_56_39), .reg_activation(reg_activation_57_39), .reg_weight(reg_weight_57_39), .reg_partial_sum(reg_psum_57_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_40( .activation_in(reg_activation_57_39), .weight_in(reg_weight_56_40), .partial_sum_in(reg_psum_56_40), .reg_activation(reg_activation_57_40), .reg_weight(reg_weight_57_40), .reg_partial_sum(reg_psum_57_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_41( .activation_in(reg_activation_57_40), .weight_in(reg_weight_56_41), .partial_sum_in(reg_psum_56_41), .reg_activation(reg_activation_57_41), .reg_weight(reg_weight_57_41), .reg_partial_sum(reg_psum_57_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_42( .activation_in(reg_activation_57_41), .weight_in(reg_weight_56_42), .partial_sum_in(reg_psum_56_42), .reg_activation(reg_activation_57_42), .reg_weight(reg_weight_57_42), .reg_partial_sum(reg_psum_57_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_43( .activation_in(reg_activation_57_42), .weight_in(reg_weight_56_43), .partial_sum_in(reg_psum_56_43), .reg_activation(reg_activation_57_43), .reg_weight(reg_weight_57_43), .reg_partial_sum(reg_psum_57_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_44( .activation_in(reg_activation_57_43), .weight_in(reg_weight_56_44), .partial_sum_in(reg_psum_56_44), .reg_activation(reg_activation_57_44), .reg_weight(reg_weight_57_44), .reg_partial_sum(reg_psum_57_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_45( .activation_in(reg_activation_57_44), .weight_in(reg_weight_56_45), .partial_sum_in(reg_psum_56_45), .reg_activation(reg_activation_57_45), .reg_weight(reg_weight_57_45), .reg_partial_sum(reg_psum_57_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_46( .activation_in(reg_activation_57_45), .weight_in(reg_weight_56_46), .partial_sum_in(reg_psum_56_46), .reg_activation(reg_activation_57_46), .reg_weight(reg_weight_57_46), .reg_partial_sum(reg_psum_57_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_47( .activation_in(reg_activation_57_46), .weight_in(reg_weight_56_47), .partial_sum_in(reg_psum_56_47), .reg_activation(reg_activation_57_47), .reg_weight(reg_weight_57_47), .reg_partial_sum(reg_psum_57_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_48( .activation_in(reg_activation_57_47), .weight_in(reg_weight_56_48), .partial_sum_in(reg_psum_56_48), .reg_activation(reg_activation_57_48), .reg_weight(reg_weight_57_48), .reg_partial_sum(reg_psum_57_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_49( .activation_in(reg_activation_57_48), .weight_in(reg_weight_56_49), .partial_sum_in(reg_psum_56_49), .reg_activation(reg_activation_57_49), .reg_weight(reg_weight_57_49), .reg_partial_sum(reg_psum_57_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_50( .activation_in(reg_activation_57_49), .weight_in(reg_weight_56_50), .partial_sum_in(reg_psum_56_50), .reg_activation(reg_activation_57_50), .reg_weight(reg_weight_57_50), .reg_partial_sum(reg_psum_57_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_51( .activation_in(reg_activation_57_50), .weight_in(reg_weight_56_51), .partial_sum_in(reg_psum_56_51), .reg_activation(reg_activation_57_51), .reg_weight(reg_weight_57_51), .reg_partial_sum(reg_psum_57_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_52( .activation_in(reg_activation_57_51), .weight_in(reg_weight_56_52), .partial_sum_in(reg_psum_56_52), .reg_activation(reg_activation_57_52), .reg_weight(reg_weight_57_52), .reg_partial_sum(reg_psum_57_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_53( .activation_in(reg_activation_57_52), .weight_in(reg_weight_56_53), .partial_sum_in(reg_psum_56_53), .reg_activation(reg_activation_57_53), .reg_weight(reg_weight_57_53), .reg_partial_sum(reg_psum_57_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_54( .activation_in(reg_activation_57_53), .weight_in(reg_weight_56_54), .partial_sum_in(reg_psum_56_54), .reg_activation(reg_activation_57_54), .reg_weight(reg_weight_57_54), .reg_partial_sum(reg_psum_57_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_55( .activation_in(reg_activation_57_54), .weight_in(reg_weight_56_55), .partial_sum_in(reg_psum_56_55), .reg_activation(reg_activation_57_55), .reg_weight(reg_weight_57_55), .reg_partial_sum(reg_psum_57_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_56( .activation_in(reg_activation_57_55), .weight_in(reg_weight_56_56), .partial_sum_in(reg_psum_56_56), .reg_activation(reg_activation_57_56), .reg_weight(reg_weight_57_56), .reg_partial_sum(reg_psum_57_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_57( .activation_in(reg_activation_57_56), .weight_in(reg_weight_56_57), .partial_sum_in(reg_psum_56_57), .reg_activation(reg_activation_57_57), .reg_weight(reg_weight_57_57), .reg_partial_sum(reg_psum_57_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_58( .activation_in(reg_activation_57_57), .weight_in(reg_weight_56_58), .partial_sum_in(reg_psum_56_58), .reg_activation(reg_activation_57_58), .reg_weight(reg_weight_57_58), .reg_partial_sum(reg_psum_57_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_59( .activation_in(reg_activation_57_58), .weight_in(reg_weight_56_59), .partial_sum_in(reg_psum_56_59), .reg_activation(reg_activation_57_59), .reg_weight(reg_weight_57_59), .reg_partial_sum(reg_psum_57_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_60( .activation_in(reg_activation_57_59), .weight_in(reg_weight_56_60), .partial_sum_in(reg_psum_56_60), .reg_activation(reg_activation_57_60), .reg_weight(reg_weight_57_60), .reg_partial_sum(reg_psum_57_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_61( .activation_in(reg_activation_57_60), .weight_in(reg_weight_56_61), .partial_sum_in(reg_psum_56_61), .reg_activation(reg_activation_57_61), .reg_weight(reg_weight_57_61), .reg_partial_sum(reg_psum_57_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_62( .activation_in(reg_activation_57_61), .weight_in(reg_weight_56_62), .partial_sum_in(reg_psum_56_62), .reg_activation(reg_activation_57_62), .reg_weight(reg_weight_57_62), .reg_partial_sum(reg_psum_57_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U57_63( .activation_in(reg_activation_57_62), .weight_in(reg_weight_56_63), .partial_sum_in(reg_psum_56_63), .reg_weight(reg_weight_57_63), .reg_partial_sum(reg_psum_57_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_0( .activation_in(in_activation_58), .weight_in(reg_weight_57_0), .partial_sum_in(reg_psum_57_0), .reg_activation(reg_activation_58_0), .reg_weight(reg_weight_58_0), .reg_partial_sum(reg_psum_58_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_1( .activation_in(reg_activation_58_0), .weight_in(reg_weight_57_1), .partial_sum_in(reg_psum_57_1), .reg_activation(reg_activation_58_1), .reg_weight(reg_weight_58_1), .reg_partial_sum(reg_psum_58_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_2( .activation_in(reg_activation_58_1), .weight_in(reg_weight_57_2), .partial_sum_in(reg_psum_57_2), .reg_activation(reg_activation_58_2), .reg_weight(reg_weight_58_2), .reg_partial_sum(reg_psum_58_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_3( .activation_in(reg_activation_58_2), .weight_in(reg_weight_57_3), .partial_sum_in(reg_psum_57_3), .reg_activation(reg_activation_58_3), .reg_weight(reg_weight_58_3), .reg_partial_sum(reg_psum_58_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_4( .activation_in(reg_activation_58_3), .weight_in(reg_weight_57_4), .partial_sum_in(reg_psum_57_4), .reg_activation(reg_activation_58_4), .reg_weight(reg_weight_58_4), .reg_partial_sum(reg_psum_58_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_5( .activation_in(reg_activation_58_4), .weight_in(reg_weight_57_5), .partial_sum_in(reg_psum_57_5), .reg_activation(reg_activation_58_5), .reg_weight(reg_weight_58_5), .reg_partial_sum(reg_psum_58_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_6( .activation_in(reg_activation_58_5), .weight_in(reg_weight_57_6), .partial_sum_in(reg_psum_57_6), .reg_activation(reg_activation_58_6), .reg_weight(reg_weight_58_6), .reg_partial_sum(reg_psum_58_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_7( .activation_in(reg_activation_58_6), .weight_in(reg_weight_57_7), .partial_sum_in(reg_psum_57_7), .reg_activation(reg_activation_58_7), .reg_weight(reg_weight_58_7), .reg_partial_sum(reg_psum_58_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_8( .activation_in(reg_activation_58_7), .weight_in(reg_weight_57_8), .partial_sum_in(reg_psum_57_8), .reg_activation(reg_activation_58_8), .reg_weight(reg_weight_58_8), .reg_partial_sum(reg_psum_58_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_9( .activation_in(reg_activation_58_8), .weight_in(reg_weight_57_9), .partial_sum_in(reg_psum_57_9), .reg_activation(reg_activation_58_9), .reg_weight(reg_weight_58_9), .reg_partial_sum(reg_psum_58_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_10( .activation_in(reg_activation_58_9), .weight_in(reg_weight_57_10), .partial_sum_in(reg_psum_57_10), .reg_activation(reg_activation_58_10), .reg_weight(reg_weight_58_10), .reg_partial_sum(reg_psum_58_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_11( .activation_in(reg_activation_58_10), .weight_in(reg_weight_57_11), .partial_sum_in(reg_psum_57_11), .reg_activation(reg_activation_58_11), .reg_weight(reg_weight_58_11), .reg_partial_sum(reg_psum_58_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_12( .activation_in(reg_activation_58_11), .weight_in(reg_weight_57_12), .partial_sum_in(reg_psum_57_12), .reg_activation(reg_activation_58_12), .reg_weight(reg_weight_58_12), .reg_partial_sum(reg_psum_58_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_13( .activation_in(reg_activation_58_12), .weight_in(reg_weight_57_13), .partial_sum_in(reg_psum_57_13), .reg_activation(reg_activation_58_13), .reg_weight(reg_weight_58_13), .reg_partial_sum(reg_psum_58_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_14( .activation_in(reg_activation_58_13), .weight_in(reg_weight_57_14), .partial_sum_in(reg_psum_57_14), .reg_activation(reg_activation_58_14), .reg_weight(reg_weight_58_14), .reg_partial_sum(reg_psum_58_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_15( .activation_in(reg_activation_58_14), .weight_in(reg_weight_57_15), .partial_sum_in(reg_psum_57_15), .reg_activation(reg_activation_58_15), .reg_weight(reg_weight_58_15), .reg_partial_sum(reg_psum_58_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_16( .activation_in(reg_activation_58_15), .weight_in(reg_weight_57_16), .partial_sum_in(reg_psum_57_16), .reg_activation(reg_activation_58_16), .reg_weight(reg_weight_58_16), .reg_partial_sum(reg_psum_58_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_17( .activation_in(reg_activation_58_16), .weight_in(reg_weight_57_17), .partial_sum_in(reg_psum_57_17), .reg_activation(reg_activation_58_17), .reg_weight(reg_weight_58_17), .reg_partial_sum(reg_psum_58_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_18( .activation_in(reg_activation_58_17), .weight_in(reg_weight_57_18), .partial_sum_in(reg_psum_57_18), .reg_activation(reg_activation_58_18), .reg_weight(reg_weight_58_18), .reg_partial_sum(reg_psum_58_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_19( .activation_in(reg_activation_58_18), .weight_in(reg_weight_57_19), .partial_sum_in(reg_psum_57_19), .reg_activation(reg_activation_58_19), .reg_weight(reg_weight_58_19), .reg_partial_sum(reg_psum_58_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_20( .activation_in(reg_activation_58_19), .weight_in(reg_weight_57_20), .partial_sum_in(reg_psum_57_20), .reg_activation(reg_activation_58_20), .reg_weight(reg_weight_58_20), .reg_partial_sum(reg_psum_58_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_21( .activation_in(reg_activation_58_20), .weight_in(reg_weight_57_21), .partial_sum_in(reg_psum_57_21), .reg_activation(reg_activation_58_21), .reg_weight(reg_weight_58_21), .reg_partial_sum(reg_psum_58_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_22( .activation_in(reg_activation_58_21), .weight_in(reg_weight_57_22), .partial_sum_in(reg_psum_57_22), .reg_activation(reg_activation_58_22), .reg_weight(reg_weight_58_22), .reg_partial_sum(reg_psum_58_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_23( .activation_in(reg_activation_58_22), .weight_in(reg_weight_57_23), .partial_sum_in(reg_psum_57_23), .reg_activation(reg_activation_58_23), .reg_weight(reg_weight_58_23), .reg_partial_sum(reg_psum_58_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_24( .activation_in(reg_activation_58_23), .weight_in(reg_weight_57_24), .partial_sum_in(reg_psum_57_24), .reg_activation(reg_activation_58_24), .reg_weight(reg_weight_58_24), .reg_partial_sum(reg_psum_58_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_25( .activation_in(reg_activation_58_24), .weight_in(reg_weight_57_25), .partial_sum_in(reg_psum_57_25), .reg_activation(reg_activation_58_25), .reg_weight(reg_weight_58_25), .reg_partial_sum(reg_psum_58_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_26( .activation_in(reg_activation_58_25), .weight_in(reg_weight_57_26), .partial_sum_in(reg_psum_57_26), .reg_activation(reg_activation_58_26), .reg_weight(reg_weight_58_26), .reg_partial_sum(reg_psum_58_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_27( .activation_in(reg_activation_58_26), .weight_in(reg_weight_57_27), .partial_sum_in(reg_psum_57_27), .reg_activation(reg_activation_58_27), .reg_weight(reg_weight_58_27), .reg_partial_sum(reg_psum_58_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_28( .activation_in(reg_activation_58_27), .weight_in(reg_weight_57_28), .partial_sum_in(reg_psum_57_28), .reg_activation(reg_activation_58_28), .reg_weight(reg_weight_58_28), .reg_partial_sum(reg_psum_58_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_29( .activation_in(reg_activation_58_28), .weight_in(reg_weight_57_29), .partial_sum_in(reg_psum_57_29), .reg_activation(reg_activation_58_29), .reg_weight(reg_weight_58_29), .reg_partial_sum(reg_psum_58_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_30( .activation_in(reg_activation_58_29), .weight_in(reg_weight_57_30), .partial_sum_in(reg_psum_57_30), .reg_activation(reg_activation_58_30), .reg_weight(reg_weight_58_30), .reg_partial_sum(reg_psum_58_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_31( .activation_in(reg_activation_58_30), .weight_in(reg_weight_57_31), .partial_sum_in(reg_psum_57_31), .reg_activation(reg_activation_58_31), .reg_weight(reg_weight_58_31), .reg_partial_sum(reg_psum_58_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_32( .activation_in(reg_activation_58_31), .weight_in(reg_weight_57_32), .partial_sum_in(reg_psum_57_32), .reg_activation(reg_activation_58_32), .reg_weight(reg_weight_58_32), .reg_partial_sum(reg_psum_58_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_33( .activation_in(reg_activation_58_32), .weight_in(reg_weight_57_33), .partial_sum_in(reg_psum_57_33), .reg_activation(reg_activation_58_33), .reg_weight(reg_weight_58_33), .reg_partial_sum(reg_psum_58_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_34( .activation_in(reg_activation_58_33), .weight_in(reg_weight_57_34), .partial_sum_in(reg_psum_57_34), .reg_activation(reg_activation_58_34), .reg_weight(reg_weight_58_34), .reg_partial_sum(reg_psum_58_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_35( .activation_in(reg_activation_58_34), .weight_in(reg_weight_57_35), .partial_sum_in(reg_psum_57_35), .reg_activation(reg_activation_58_35), .reg_weight(reg_weight_58_35), .reg_partial_sum(reg_psum_58_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_36( .activation_in(reg_activation_58_35), .weight_in(reg_weight_57_36), .partial_sum_in(reg_psum_57_36), .reg_activation(reg_activation_58_36), .reg_weight(reg_weight_58_36), .reg_partial_sum(reg_psum_58_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_37( .activation_in(reg_activation_58_36), .weight_in(reg_weight_57_37), .partial_sum_in(reg_psum_57_37), .reg_activation(reg_activation_58_37), .reg_weight(reg_weight_58_37), .reg_partial_sum(reg_psum_58_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_38( .activation_in(reg_activation_58_37), .weight_in(reg_weight_57_38), .partial_sum_in(reg_psum_57_38), .reg_activation(reg_activation_58_38), .reg_weight(reg_weight_58_38), .reg_partial_sum(reg_psum_58_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_39( .activation_in(reg_activation_58_38), .weight_in(reg_weight_57_39), .partial_sum_in(reg_psum_57_39), .reg_activation(reg_activation_58_39), .reg_weight(reg_weight_58_39), .reg_partial_sum(reg_psum_58_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_40( .activation_in(reg_activation_58_39), .weight_in(reg_weight_57_40), .partial_sum_in(reg_psum_57_40), .reg_activation(reg_activation_58_40), .reg_weight(reg_weight_58_40), .reg_partial_sum(reg_psum_58_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_41( .activation_in(reg_activation_58_40), .weight_in(reg_weight_57_41), .partial_sum_in(reg_psum_57_41), .reg_activation(reg_activation_58_41), .reg_weight(reg_weight_58_41), .reg_partial_sum(reg_psum_58_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_42( .activation_in(reg_activation_58_41), .weight_in(reg_weight_57_42), .partial_sum_in(reg_psum_57_42), .reg_activation(reg_activation_58_42), .reg_weight(reg_weight_58_42), .reg_partial_sum(reg_psum_58_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_43( .activation_in(reg_activation_58_42), .weight_in(reg_weight_57_43), .partial_sum_in(reg_psum_57_43), .reg_activation(reg_activation_58_43), .reg_weight(reg_weight_58_43), .reg_partial_sum(reg_psum_58_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_44( .activation_in(reg_activation_58_43), .weight_in(reg_weight_57_44), .partial_sum_in(reg_psum_57_44), .reg_activation(reg_activation_58_44), .reg_weight(reg_weight_58_44), .reg_partial_sum(reg_psum_58_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_45( .activation_in(reg_activation_58_44), .weight_in(reg_weight_57_45), .partial_sum_in(reg_psum_57_45), .reg_activation(reg_activation_58_45), .reg_weight(reg_weight_58_45), .reg_partial_sum(reg_psum_58_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_46( .activation_in(reg_activation_58_45), .weight_in(reg_weight_57_46), .partial_sum_in(reg_psum_57_46), .reg_activation(reg_activation_58_46), .reg_weight(reg_weight_58_46), .reg_partial_sum(reg_psum_58_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_47( .activation_in(reg_activation_58_46), .weight_in(reg_weight_57_47), .partial_sum_in(reg_psum_57_47), .reg_activation(reg_activation_58_47), .reg_weight(reg_weight_58_47), .reg_partial_sum(reg_psum_58_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_48( .activation_in(reg_activation_58_47), .weight_in(reg_weight_57_48), .partial_sum_in(reg_psum_57_48), .reg_activation(reg_activation_58_48), .reg_weight(reg_weight_58_48), .reg_partial_sum(reg_psum_58_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_49( .activation_in(reg_activation_58_48), .weight_in(reg_weight_57_49), .partial_sum_in(reg_psum_57_49), .reg_activation(reg_activation_58_49), .reg_weight(reg_weight_58_49), .reg_partial_sum(reg_psum_58_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_50( .activation_in(reg_activation_58_49), .weight_in(reg_weight_57_50), .partial_sum_in(reg_psum_57_50), .reg_activation(reg_activation_58_50), .reg_weight(reg_weight_58_50), .reg_partial_sum(reg_psum_58_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_51( .activation_in(reg_activation_58_50), .weight_in(reg_weight_57_51), .partial_sum_in(reg_psum_57_51), .reg_activation(reg_activation_58_51), .reg_weight(reg_weight_58_51), .reg_partial_sum(reg_psum_58_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_52( .activation_in(reg_activation_58_51), .weight_in(reg_weight_57_52), .partial_sum_in(reg_psum_57_52), .reg_activation(reg_activation_58_52), .reg_weight(reg_weight_58_52), .reg_partial_sum(reg_psum_58_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_53( .activation_in(reg_activation_58_52), .weight_in(reg_weight_57_53), .partial_sum_in(reg_psum_57_53), .reg_activation(reg_activation_58_53), .reg_weight(reg_weight_58_53), .reg_partial_sum(reg_psum_58_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_54( .activation_in(reg_activation_58_53), .weight_in(reg_weight_57_54), .partial_sum_in(reg_psum_57_54), .reg_activation(reg_activation_58_54), .reg_weight(reg_weight_58_54), .reg_partial_sum(reg_psum_58_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_55( .activation_in(reg_activation_58_54), .weight_in(reg_weight_57_55), .partial_sum_in(reg_psum_57_55), .reg_activation(reg_activation_58_55), .reg_weight(reg_weight_58_55), .reg_partial_sum(reg_psum_58_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_56( .activation_in(reg_activation_58_55), .weight_in(reg_weight_57_56), .partial_sum_in(reg_psum_57_56), .reg_activation(reg_activation_58_56), .reg_weight(reg_weight_58_56), .reg_partial_sum(reg_psum_58_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_57( .activation_in(reg_activation_58_56), .weight_in(reg_weight_57_57), .partial_sum_in(reg_psum_57_57), .reg_activation(reg_activation_58_57), .reg_weight(reg_weight_58_57), .reg_partial_sum(reg_psum_58_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_58( .activation_in(reg_activation_58_57), .weight_in(reg_weight_57_58), .partial_sum_in(reg_psum_57_58), .reg_activation(reg_activation_58_58), .reg_weight(reg_weight_58_58), .reg_partial_sum(reg_psum_58_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_59( .activation_in(reg_activation_58_58), .weight_in(reg_weight_57_59), .partial_sum_in(reg_psum_57_59), .reg_activation(reg_activation_58_59), .reg_weight(reg_weight_58_59), .reg_partial_sum(reg_psum_58_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_60( .activation_in(reg_activation_58_59), .weight_in(reg_weight_57_60), .partial_sum_in(reg_psum_57_60), .reg_activation(reg_activation_58_60), .reg_weight(reg_weight_58_60), .reg_partial_sum(reg_psum_58_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_61( .activation_in(reg_activation_58_60), .weight_in(reg_weight_57_61), .partial_sum_in(reg_psum_57_61), .reg_activation(reg_activation_58_61), .reg_weight(reg_weight_58_61), .reg_partial_sum(reg_psum_58_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_62( .activation_in(reg_activation_58_61), .weight_in(reg_weight_57_62), .partial_sum_in(reg_psum_57_62), .reg_activation(reg_activation_58_62), .reg_weight(reg_weight_58_62), .reg_partial_sum(reg_psum_58_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U58_63( .activation_in(reg_activation_58_62), .weight_in(reg_weight_57_63), .partial_sum_in(reg_psum_57_63), .reg_weight(reg_weight_58_63), .reg_partial_sum(reg_psum_58_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_0( .activation_in(in_activation_59), .weight_in(reg_weight_58_0), .partial_sum_in(reg_psum_58_0), .reg_activation(reg_activation_59_0), .reg_weight(reg_weight_59_0), .reg_partial_sum(reg_psum_59_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_1( .activation_in(reg_activation_59_0), .weight_in(reg_weight_58_1), .partial_sum_in(reg_psum_58_1), .reg_activation(reg_activation_59_1), .reg_weight(reg_weight_59_1), .reg_partial_sum(reg_psum_59_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_2( .activation_in(reg_activation_59_1), .weight_in(reg_weight_58_2), .partial_sum_in(reg_psum_58_2), .reg_activation(reg_activation_59_2), .reg_weight(reg_weight_59_2), .reg_partial_sum(reg_psum_59_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_3( .activation_in(reg_activation_59_2), .weight_in(reg_weight_58_3), .partial_sum_in(reg_psum_58_3), .reg_activation(reg_activation_59_3), .reg_weight(reg_weight_59_3), .reg_partial_sum(reg_psum_59_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_4( .activation_in(reg_activation_59_3), .weight_in(reg_weight_58_4), .partial_sum_in(reg_psum_58_4), .reg_activation(reg_activation_59_4), .reg_weight(reg_weight_59_4), .reg_partial_sum(reg_psum_59_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_5( .activation_in(reg_activation_59_4), .weight_in(reg_weight_58_5), .partial_sum_in(reg_psum_58_5), .reg_activation(reg_activation_59_5), .reg_weight(reg_weight_59_5), .reg_partial_sum(reg_psum_59_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_6( .activation_in(reg_activation_59_5), .weight_in(reg_weight_58_6), .partial_sum_in(reg_psum_58_6), .reg_activation(reg_activation_59_6), .reg_weight(reg_weight_59_6), .reg_partial_sum(reg_psum_59_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_7( .activation_in(reg_activation_59_6), .weight_in(reg_weight_58_7), .partial_sum_in(reg_psum_58_7), .reg_activation(reg_activation_59_7), .reg_weight(reg_weight_59_7), .reg_partial_sum(reg_psum_59_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_8( .activation_in(reg_activation_59_7), .weight_in(reg_weight_58_8), .partial_sum_in(reg_psum_58_8), .reg_activation(reg_activation_59_8), .reg_weight(reg_weight_59_8), .reg_partial_sum(reg_psum_59_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_9( .activation_in(reg_activation_59_8), .weight_in(reg_weight_58_9), .partial_sum_in(reg_psum_58_9), .reg_activation(reg_activation_59_9), .reg_weight(reg_weight_59_9), .reg_partial_sum(reg_psum_59_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_10( .activation_in(reg_activation_59_9), .weight_in(reg_weight_58_10), .partial_sum_in(reg_psum_58_10), .reg_activation(reg_activation_59_10), .reg_weight(reg_weight_59_10), .reg_partial_sum(reg_psum_59_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_11( .activation_in(reg_activation_59_10), .weight_in(reg_weight_58_11), .partial_sum_in(reg_psum_58_11), .reg_activation(reg_activation_59_11), .reg_weight(reg_weight_59_11), .reg_partial_sum(reg_psum_59_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_12( .activation_in(reg_activation_59_11), .weight_in(reg_weight_58_12), .partial_sum_in(reg_psum_58_12), .reg_activation(reg_activation_59_12), .reg_weight(reg_weight_59_12), .reg_partial_sum(reg_psum_59_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_13( .activation_in(reg_activation_59_12), .weight_in(reg_weight_58_13), .partial_sum_in(reg_psum_58_13), .reg_activation(reg_activation_59_13), .reg_weight(reg_weight_59_13), .reg_partial_sum(reg_psum_59_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_14( .activation_in(reg_activation_59_13), .weight_in(reg_weight_58_14), .partial_sum_in(reg_psum_58_14), .reg_activation(reg_activation_59_14), .reg_weight(reg_weight_59_14), .reg_partial_sum(reg_psum_59_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_15( .activation_in(reg_activation_59_14), .weight_in(reg_weight_58_15), .partial_sum_in(reg_psum_58_15), .reg_activation(reg_activation_59_15), .reg_weight(reg_weight_59_15), .reg_partial_sum(reg_psum_59_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_16( .activation_in(reg_activation_59_15), .weight_in(reg_weight_58_16), .partial_sum_in(reg_psum_58_16), .reg_activation(reg_activation_59_16), .reg_weight(reg_weight_59_16), .reg_partial_sum(reg_psum_59_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_17( .activation_in(reg_activation_59_16), .weight_in(reg_weight_58_17), .partial_sum_in(reg_psum_58_17), .reg_activation(reg_activation_59_17), .reg_weight(reg_weight_59_17), .reg_partial_sum(reg_psum_59_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_18( .activation_in(reg_activation_59_17), .weight_in(reg_weight_58_18), .partial_sum_in(reg_psum_58_18), .reg_activation(reg_activation_59_18), .reg_weight(reg_weight_59_18), .reg_partial_sum(reg_psum_59_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_19( .activation_in(reg_activation_59_18), .weight_in(reg_weight_58_19), .partial_sum_in(reg_psum_58_19), .reg_activation(reg_activation_59_19), .reg_weight(reg_weight_59_19), .reg_partial_sum(reg_psum_59_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_20( .activation_in(reg_activation_59_19), .weight_in(reg_weight_58_20), .partial_sum_in(reg_psum_58_20), .reg_activation(reg_activation_59_20), .reg_weight(reg_weight_59_20), .reg_partial_sum(reg_psum_59_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_21( .activation_in(reg_activation_59_20), .weight_in(reg_weight_58_21), .partial_sum_in(reg_psum_58_21), .reg_activation(reg_activation_59_21), .reg_weight(reg_weight_59_21), .reg_partial_sum(reg_psum_59_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_22( .activation_in(reg_activation_59_21), .weight_in(reg_weight_58_22), .partial_sum_in(reg_psum_58_22), .reg_activation(reg_activation_59_22), .reg_weight(reg_weight_59_22), .reg_partial_sum(reg_psum_59_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_23( .activation_in(reg_activation_59_22), .weight_in(reg_weight_58_23), .partial_sum_in(reg_psum_58_23), .reg_activation(reg_activation_59_23), .reg_weight(reg_weight_59_23), .reg_partial_sum(reg_psum_59_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_24( .activation_in(reg_activation_59_23), .weight_in(reg_weight_58_24), .partial_sum_in(reg_psum_58_24), .reg_activation(reg_activation_59_24), .reg_weight(reg_weight_59_24), .reg_partial_sum(reg_psum_59_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_25( .activation_in(reg_activation_59_24), .weight_in(reg_weight_58_25), .partial_sum_in(reg_psum_58_25), .reg_activation(reg_activation_59_25), .reg_weight(reg_weight_59_25), .reg_partial_sum(reg_psum_59_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_26( .activation_in(reg_activation_59_25), .weight_in(reg_weight_58_26), .partial_sum_in(reg_psum_58_26), .reg_activation(reg_activation_59_26), .reg_weight(reg_weight_59_26), .reg_partial_sum(reg_psum_59_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_27( .activation_in(reg_activation_59_26), .weight_in(reg_weight_58_27), .partial_sum_in(reg_psum_58_27), .reg_activation(reg_activation_59_27), .reg_weight(reg_weight_59_27), .reg_partial_sum(reg_psum_59_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_28( .activation_in(reg_activation_59_27), .weight_in(reg_weight_58_28), .partial_sum_in(reg_psum_58_28), .reg_activation(reg_activation_59_28), .reg_weight(reg_weight_59_28), .reg_partial_sum(reg_psum_59_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_29( .activation_in(reg_activation_59_28), .weight_in(reg_weight_58_29), .partial_sum_in(reg_psum_58_29), .reg_activation(reg_activation_59_29), .reg_weight(reg_weight_59_29), .reg_partial_sum(reg_psum_59_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_30( .activation_in(reg_activation_59_29), .weight_in(reg_weight_58_30), .partial_sum_in(reg_psum_58_30), .reg_activation(reg_activation_59_30), .reg_weight(reg_weight_59_30), .reg_partial_sum(reg_psum_59_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_31( .activation_in(reg_activation_59_30), .weight_in(reg_weight_58_31), .partial_sum_in(reg_psum_58_31), .reg_activation(reg_activation_59_31), .reg_weight(reg_weight_59_31), .reg_partial_sum(reg_psum_59_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_32( .activation_in(reg_activation_59_31), .weight_in(reg_weight_58_32), .partial_sum_in(reg_psum_58_32), .reg_activation(reg_activation_59_32), .reg_weight(reg_weight_59_32), .reg_partial_sum(reg_psum_59_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_33( .activation_in(reg_activation_59_32), .weight_in(reg_weight_58_33), .partial_sum_in(reg_psum_58_33), .reg_activation(reg_activation_59_33), .reg_weight(reg_weight_59_33), .reg_partial_sum(reg_psum_59_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_34( .activation_in(reg_activation_59_33), .weight_in(reg_weight_58_34), .partial_sum_in(reg_psum_58_34), .reg_activation(reg_activation_59_34), .reg_weight(reg_weight_59_34), .reg_partial_sum(reg_psum_59_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_35( .activation_in(reg_activation_59_34), .weight_in(reg_weight_58_35), .partial_sum_in(reg_psum_58_35), .reg_activation(reg_activation_59_35), .reg_weight(reg_weight_59_35), .reg_partial_sum(reg_psum_59_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_36( .activation_in(reg_activation_59_35), .weight_in(reg_weight_58_36), .partial_sum_in(reg_psum_58_36), .reg_activation(reg_activation_59_36), .reg_weight(reg_weight_59_36), .reg_partial_sum(reg_psum_59_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_37( .activation_in(reg_activation_59_36), .weight_in(reg_weight_58_37), .partial_sum_in(reg_psum_58_37), .reg_activation(reg_activation_59_37), .reg_weight(reg_weight_59_37), .reg_partial_sum(reg_psum_59_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_38( .activation_in(reg_activation_59_37), .weight_in(reg_weight_58_38), .partial_sum_in(reg_psum_58_38), .reg_activation(reg_activation_59_38), .reg_weight(reg_weight_59_38), .reg_partial_sum(reg_psum_59_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_39( .activation_in(reg_activation_59_38), .weight_in(reg_weight_58_39), .partial_sum_in(reg_psum_58_39), .reg_activation(reg_activation_59_39), .reg_weight(reg_weight_59_39), .reg_partial_sum(reg_psum_59_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_40( .activation_in(reg_activation_59_39), .weight_in(reg_weight_58_40), .partial_sum_in(reg_psum_58_40), .reg_activation(reg_activation_59_40), .reg_weight(reg_weight_59_40), .reg_partial_sum(reg_psum_59_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_41( .activation_in(reg_activation_59_40), .weight_in(reg_weight_58_41), .partial_sum_in(reg_psum_58_41), .reg_activation(reg_activation_59_41), .reg_weight(reg_weight_59_41), .reg_partial_sum(reg_psum_59_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_42( .activation_in(reg_activation_59_41), .weight_in(reg_weight_58_42), .partial_sum_in(reg_psum_58_42), .reg_activation(reg_activation_59_42), .reg_weight(reg_weight_59_42), .reg_partial_sum(reg_psum_59_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_43( .activation_in(reg_activation_59_42), .weight_in(reg_weight_58_43), .partial_sum_in(reg_psum_58_43), .reg_activation(reg_activation_59_43), .reg_weight(reg_weight_59_43), .reg_partial_sum(reg_psum_59_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_44( .activation_in(reg_activation_59_43), .weight_in(reg_weight_58_44), .partial_sum_in(reg_psum_58_44), .reg_activation(reg_activation_59_44), .reg_weight(reg_weight_59_44), .reg_partial_sum(reg_psum_59_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_45( .activation_in(reg_activation_59_44), .weight_in(reg_weight_58_45), .partial_sum_in(reg_psum_58_45), .reg_activation(reg_activation_59_45), .reg_weight(reg_weight_59_45), .reg_partial_sum(reg_psum_59_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_46( .activation_in(reg_activation_59_45), .weight_in(reg_weight_58_46), .partial_sum_in(reg_psum_58_46), .reg_activation(reg_activation_59_46), .reg_weight(reg_weight_59_46), .reg_partial_sum(reg_psum_59_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_47( .activation_in(reg_activation_59_46), .weight_in(reg_weight_58_47), .partial_sum_in(reg_psum_58_47), .reg_activation(reg_activation_59_47), .reg_weight(reg_weight_59_47), .reg_partial_sum(reg_psum_59_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_48( .activation_in(reg_activation_59_47), .weight_in(reg_weight_58_48), .partial_sum_in(reg_psum_58_48), .reg_activation(reg_activation_59_48), .reg_weight(reg_weight_59_48), .reg_partial_sum(reg_psum_59_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_49( .activation_in(reg_activation_59_48), .weight_in(reg_weight_58_49), .partial_sum_in(reg_psum_58_49), .reg_activation(reg_activation_59_49), .reg_weight(reg_weight_59_49), .reg_partial_sum(reg_psum_59_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_50( .activation_in(reg_activation_59_49), .weight_in(reg_weight_58_50), .partial_sum_in(reg_psum_58_50), .reg_activation(reg_activation_59_50), .reg_weight(reg_weight_59_50), .reg_partial_sum(reg_psum_59_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_51( .activation_in(reg_activation_59_50), .weight_in(reg_weight_58_51), .partial_sum_in(reg_psum_58_51), .reg_activation(reg_activation_59_51), .reg_weight(reg_weight_59_51), .reg_partial_sum(reg_psum_59_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_52( .activation_in(reg_activation_59_51), .weight_in(reg_weight_58_52), .partial_sum_in(reg_psum_58_52), .reg_activation(reg_activation_59_52), .reg_weight(reg_weight_59_52), .reg_partial_sum(reg_psum_59_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_53( .activation_in(reg_activation_59_52), .weight_in(reg_weight_58_53), .partial_sum_in(reg_psum_58_53), .reg_activation(reg_activation_59_53), .reg_weight(reg_weight_59_53), .reg_partial_sum(reg_psum_59_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_54( .activation_in(reg_activation_59_53), .weight_in(reg_weight_58_54), .partial_sum_in(reg_psum_58_54), .reg_activation(reg_activation_59_54), .reg_weight(reg_weight_59_54), .reg_partial_sum(reg_psum_59_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_55( .activation_in(reg_activation_59_54), .weight_in(reg_weight_58_55), .partial_sum_in(reg_psum_58_55), .reg_activation(reg_activation_59_55), .reg_weight(reg_weight_59_55), .reg_partial_sum(reg_psum_59_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_56( .activation_in(reg_activation_59_55), .weight_in(reg_weight_58_56), .partial_sum_in(reg_psum_58_56), .reg_activation(reg_activation_59_56), .reg_weight(reg_weight_59_56), .reg_partial_sum(reg_psum_59_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_57( .activation_in(reg_activation_59_56), .weight_in(reg_weight_58_57), .partial_sum_in(reg_psum_58_57), .reg_activation(reg_activation_59_57), .reg_weight(reg_weight_59_57), .reg_partial_sum(reg_psum_59_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_58( .activation_in(reg_activation_59_57), .weight_in(reg_weight_58_58), .partial_sum_in(reg_psum_58_58), .reg_activation(reg_activation_59_58), .reg_weight(reg_weight_59_58), .reg_partial_sum(reg_psum_59_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_59( .activation_in(reg_activation_59_58), .weight_in(reg_weight_58_59), .partial_sum_in(reg_psum_58_59), .reg_activation(reg_activation_59_59), .reg_weight(reg_weight_59_59), .reg_partial_sum(reg_psum_59_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_60( .activation_in(reg_activation_59_59), .weight_in(reg_weight_58_60), .partial_sum_in(reg_psum_58_60), .reg_activation(reg_activation_59_60), .reg_weight(reg_weight_59_60), .reg_partial_sum(reg_psum_59_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_61( .activation_in(reg_activation_59_60), .weight_in(reg_weight_58_61), .partial_sum_in(reg_psum_58_61), .reg_activation(reg_activation_59_61), .reg_weight(reg_weight_59_61), .reg_partial_sum(reg_psum_59_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_62( .activation_in(reg_activation_59_61), .weight_in(reg_weight_58_62), .partial_sum_in(reg_psum_58_62), .reg_activation(reg_activation_59_62), .reg_weight(reg_weight_59_62), .reg_partial_sum(reg_psum_59_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U59_63( .activation_in(reg_activation_59_62), .weight_in(reg_weight_58_63), .partial_sum_in(reg_psum_58_63), .reg_weight(reg_weight_59_63), .reg_partial_sum(reg_psum_59_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_0( .activation_in(in_activation_60), .weight_in(reg_weight_59_0), .partial_sum_in(reg_psum_59_0), .reg_activation(reg_activation_60_0), .reg_weight(reg_weight_60_0), .reg_partial_sum(reg_psum_60_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_1( .activation_in(reg_activation_60_0), .weight_in(reg_weight_59_1), .partial_sum_in(reg_psum_59_1), .reg_activation(reg_activation_60_1), .reg_weight(reg_weight_60_1), .reg_partial_sum(reg_psum_60_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_2( .activation_in(reg_activation_60_1), .weight_in(reg_weight_59_2), .partial_sum_in(reg_psum_59_2), .reg_activation(reg_activation_60_2), .reg_weight(reg_weight_60_2), .reg_partial_sum(reg_psum_60_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_3( .activation_in(reg_activation_60_2), .weight_in(reg_weight_59_3), .partial_sum_in(reg_psum_59_3), .reg_activation(reg_activation_60_3), .reg_weight(reg_weight_60_3), .reg_partial_sum(reg_psum_60_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_4( .activation_in(reg_activation_60_3), .weight_in(reg_weight_59_4), .partial_sum_in(reg_psum_59_4), .reg_activation(reg_activation_60_4), .reg_weight(reg_weight_60_4), .reg_partial_sum(reg_psum_60_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_5( .activation_in(reg_activation_60_4), .weight_in(reg_weight_59_5), .partial_sum_in(reg_psum_59_5), .reg_activation(reg_activation_60_5), .reg_weight(reg_weight_60_5), .reg_partial_sum(reg_psum_60_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_6( .activation_in(reg_activation_60_5), .weight_in(reg_weight_59_6), .partial_sum_in(reg_psum_59_6), .reg_activation(reg_activation_60_6), .reg_weight(reg_weight_60_6), .reg_partial_sum(reg_psum_60_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_7( .activation_in(reg_activation_60_6), .weight_in(reg_weight_59_7), .partial_sum_in(reg_psum_59_7), .reg_activation(reg_activation_60_7), .reg_weight(reg_weight_60_7), .reg_partial_sum(reg_psum_60_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_8( .activation_in(reg_activation_60_7), .weight_in(reg_weight_59_8), .partial_sum_in(reg_psum_59_8), .reg_activation(reg_activation_60_8), .reg_weight(reg_weight_60_8), .reg_partial_sum(reg_psum_60_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_9( .activation_in(reg_activation_60_8), .weight_in(reg_weight_59_9), .partial_sum_in(reg_psum_59_9), .reg_activation(reg_activation_60_9), .reg_weight(reg_weight_60_9), .reg_partial_sum(reg_psum_60_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_10( .activation_in(reg_activation_60_9), .weight_in(reg_weight_59_10), .partial_sum_in(reg_psum_59_10), .reg_activation(reg_activation_60_10), .reg_weight(reg_weight_60_10), .reg_partial_sum(reg_psum_60_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_11( .activation_in(reg_activation_60_10), .weight_in(reg_weight_59_11), .partial_sum_in(reg_psum_59_11), .reg_activation(reg_activation_60_11), .reg_weight(reg_weight_60_11), .reg_partial_sum(reg_psum_60_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_12( .activation_in(reg_activation_60_11), .weight_in(reg_weight_59_12), .partial_sum_in(reg_psum_59_12), .reg_activation(reg_activation_60_12), .reg_weight(reg_weight_60_12), .reg_partial_sum(reg_psum_60_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_13( .activation_in(reg_activation_60_12), .weight_in(reg_weight_59_13), .partial_sum_in(reg_psum_59_13), .reg_activation(reg_activation_60_13), .reg_weight(reg_weight_60_13), .reg_partial_sum(reg_psum_60_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_14( .activation_in(reg_activation_60_13), .weight_in(reg_weight_59_14), .partial_sum_in(reg_psum_59_14), .reg_activation(reg_activation_60_14), .reg_weight(reg_weight_60_14), .reg_partial_sum(reg_psum_60_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_15( .activation_in(reg_activation_60_14), .weight_in(reg_weight_59_15), .partial_sum_in(reg_psum_59_15), .reg_activation(reg_activation_60_15), .reg_weight(reg_weight_60_15), .reg_partial_sum(reg_psum_60_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_16( .activation_in(reg_activation_60_15), .weight_in(reg_weight_59_16), .partial_sum_in(reg_psum_59_16), .reg_activation(reg_activation_60_16), .reg_weight(reg_weight_60_16), .reg_partial_sum(reg_psum_60_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_17( .activation_in(reg_activation_60_16), .weight_in(reg_weight_59_17), .partial_sum_in(reg_psum_59_17), .reg_activation(reg_activation_60_17), .reg_weight(reg_weight_60_17), .reg_partial_sum(reg_psum_60_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_18( .activation_in(reg_activation_60_17), .weight_in(reg_weight_59_18), .partial_sum_in(reg_psum_59_18), .reg_activation(reg_activation_60_18), .reg_weight(reg_weight_60_18), .reg_partial_sum(reg_psum_60_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_19( .activation_in(reg_activation_60_18), .weight_in(reg_weight_59_19), .partial_sum_in(reg_psum_59_19), .reg_activation(reg_activation_60_19), .reg_weight(reg_weight_60_19), .reg_partial_sum(reg_psum_60_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_20( .activation_in(reg_activation_60_19), .weight_in(reg_weight_59_20), .partial_sum_in(reg_psum_59_20), .reg_activation(reg_activation_60_20), .reg_weight(reg_weight_60_20), .reg_partial_sum(reg_psum_60_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_21( .activation_in(reg_activation_60_20), .weight_in(reg_weight_59_21), .partial_sum_in(reg_psum_59_21), .reg_activation(reg_activation_60_21), .reg_weight(reg_weight_60_21), .reg_partial_sum(reg_psum_60_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_22( .activation_in(reg_activation_60_21), .weight_in(reg_weight_59_22), .partial_sum_in(reg_psum_59_22), .reg_activation(reg_activation_60_22), .reg_weight(reg_weight_60_22), .reg_partial_sum(reg_psum_60_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_23( .activation_in(reg_activation_60_22), .weight_in(reg_weight_59_23), .partial_sum_in(reg_psum_59_23), .reg_activation(reg_activation_60_23), .reg_weight(reg_weight_60_23), .reg_partial_sum(reg_psum_60_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_24( .activation_in(reg_activation_60_23), .weight_in(reg_weight_59_24), .partial_sum_in(reg_psum_59_24), .reg_activation(reg_activation_60_24), .reg_weight(reg_weight_60_24), .reg_partial_sum(reg_psum_60_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_25( .activation_in(reg_activation_60_24), .weight_in(reg_weight_59_25), .partial_sum_in(reg_psum_59_25), .reg_activation(reg_activation_60_25), .reg_weight(reg_weight_60_25), .reg_partial_sum(reg_psum_60_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_26( .activation_in(reg_activation_60_25), .weight_in(reg_weight_59_26), .partial_sum_in(reg_psum_59_26), .reg_activation(reg_activation_60_26), .reg_weight(reg_weight_60_26), .reg_partial_sum(reg_psum_60_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_27( .activation_in(reg_activation_60_26), .weight_in(reg_weight_59_27), .partial_sum_in(reg_psum_59_27), .reg_activation(reg_activation_60_27), .reg_weight(reg_weight_60_27), .reg_partial_sum(reg_psum_60_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_28( .activation_in(reg_activation_60_27), .weight_in(reg_weight_59_28), .partial_sum_in(reg_psum_59_28), .reg_activation(reg_activation_60_28), .reg_weight(reg_weight_60_28), .reg_partial_sum(reg_psum_60_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_29( .activation_in(reg_activation_60_28), .weight_in(reg_weight_59_29), .partial_sum_in(reg_psum_59_29), .reg_activation(reg_activation_60_29), .reg_weight(reg_weight_60_29), .reg_partial_sum(reg_psum_60_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_30( .activation_in(reg_activation_60_29), .weight_in(reg_weight_59_30), .partial_sum_in(reg_psum_59_30), .reg_activation(reg_activation_60_30), .reg_weight(reg_weight_60_30), .reg_partial_sum(reg_psum_60_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_31( .activation_in(reg_activation_60_30), .weight_in(reg_weight_59_31), .partial_sum_in(reg_psum_59_31), .reg_activation(reg_activation_60_31), .reg_weight(reg_weight_60_31), .reg_partial_sum(reg_psum_60_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_32( .activation_in(reg_activation_60_31), .weight_in(reg_weight_59_32), .partial_sum_in(reg_psum_59_32), .reg_activation(reg_activation_60_32), .reg_weight(reg_weight_60_32), .reg_partial_sum(reg_psum_60_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_33( .activation_in(reg_activation_60_32), .weight_in(reg_weight_59_33), .partial_sum_in(reg_psum_59_33), .reg_activation(reg_activation_60_33), .reg_weight(reg_weight_60_33), .reg_partial_sum(reg_psum_60_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_34( .activation_in(reg_activation_60_33), .weight_in(reg_weight_59_34), .partial_sum_in(reg_psum_59_34), .reg_activation(reg_activation_60_34), .reg_weight(reg_weight_60_34), .reg_partial_sum(reg_psum_60_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_35( .activation_in(reg_activation_60_34), .weight_in(reg_weight_59_35), .partial_sum_in(reg_psum_59_35), .reg_activation(reg_activation_60_35), .reg_weight(reg_weight_60_35), .reg_partial_sum(reg_psum_60_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_36( .activation_in(reg_activation_60_35), .weight_in(reg_weight_59_36), .partial_sum_in(reg_psum_59_36), .reg_activation(reg_activation_60_36), .reg_weight(reg_weight_60_36), .reg_partial_sum(reg_psum_60_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_37( .activation_in(reg_activation_60_36), .weight_in(reg_weight_59_37), .partial_sum_in(reg_psum_59_37), .reg_activation(reg_activation_60_37), .reg_weight(reg_weight_60_37), .reg_partial_sum(reg_psum_60_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_38( .activation_in(reg_activation_60_37), .weight_in(reg_weight_59_38), .partial_sum_in(reg_psum_59_38), .reg_activation(reg_activation_60_38), .reg_weight(reg_weight_60_38), .reg_partial_sum(reg_psum_60_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_39( .activation_in(reg_activation_60_38), .weight_in(reg_weight_59_39), .partial_sum_in(reg_psum_59_39), .reg_activation(reg_activation_60_39), .reg_weight(reg_weight_60_39), .reg_partial_sum(reg_psum_60_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_40( .activation_in(reg_activation_60_39), .weight_in(reg_weight_59_40), .partial_sum_in(reg_psum_59_40), .reg_activation(reg_activation_60_40), .reg_weight(reg_weight_60_40), .reg_partial_sum(reg_psum_60_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_41( .activation_in(reg_activation_60_40), .weight_in(reg_weight_59_41), .partial_sum_in(reg_psum_59_41), .reg_activation(reg_activation_60_41), .reg_weight(reg_weight_60_41), .reg_partial_sum(reg_psum_60_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_42( .activation_in(reg_activation_60_41), .weight_in(reg_weight_59_42), .partial_sum_in(reg_psum_59_42), .reg_activation(reg_activation_60_42), .reg_weight(reg_weight_60_42), .reg_partial_sum(reg_psum_60_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_43( .activation_in(reg_activation_60_42), .weight_in(reg_weight_59_43), .partial_sum_in(reg_psum_59_43), .reg_activation(reg_activation_60_43), .reg_weight(reg_weight_60_43), .reg_partial_sum(reg_psum_60_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_44( .activation_in(reg_activation_60_43), .weight_in(reg_weight_59_44), .partial_sum_in(reg_psum_59_44), .reg_activation(reg_activation_60_44), .reg_weight(reg_weight_60_44), .reg_partial_sum(reg_psum_60_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_45( .activation_in(reg_activation_60_44), .weight_in(reg_weight_59_45), .partial_sum_in(reg_psum_59_45), .reg_activation(reg_activation_60_45), .reg_weight(reg_weight_60_45), .reg_partial_sum(reg_psum_60_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_46( .activation_in(reg_activation_60_45), .weight_in(reg_weight_59_46), .partial_sum_in(reg_psum_59_46), .reg_activation(reg_activation_60_46), .reg_weight(reg_weight_60_46), .reg_partial_sum(reg_psum_60_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_47( .activation_in(reg_activation_60_46), .weight_in(reg_weight_59_47), .partial_sum_in(reg_psum_59_47), .reg_activation(reg_activation_60_47), .reg_weight(reg_weight_60_47), .reg_partial_sum(reg_psum_60_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_48( .activation_in(reg_activation_60_47), .weight_in(reg_weight_59_48), .partial_sum_in(reg_psum_59_48), .reg_activation(reg_activation_60_48), .reg_weight(reg_weight_60_48), .reg_partial_sum(reg_psum_60_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_49( .activation_in(reg_activation_60_48), .weight_in(reg_weight_59_49), .partial_sum_in(reg_psum_59_49), .reg_activation(reg_activation_60_49), .reg_weight(reg_weight_60_49), .reg_partial_sum(reg_psum_60_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_50( .activation_in(reg_activation_60_49), .weight_in(reg_weight_59_50), .partial_sum_in(reg_psum_59_50), .reg_activation(reg_activation_60_50), .reg_weight(reg_weight_60_50), .reg_partial_sum(reg_psum_60_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_51( .activation_in(reg_activation_60_50), .weight_in(reg_weight_59_51), .partial_sum_in(reg_psum_59_51), .reg_activation(reg_activation_60_51), .reg_weight(reg_weight_60_51), .reg_partial_sum(reg_psum_60_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_52( .activation_in(reg_activation_60_51), .weight_in(reg_weight_59_52), .partial_sum_in(reg_psum_59_52), .reg_activation(reg_activation_60_52), .reg_weight(reg_weight_60_52), .reg_partial_sum(reg_psum_60_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_53( .activation_in(reg_activation_60_52), .weight_in(reg_weight_59_53), .partial_sum_in(reg_psum_59_53), .reg_activation(reg_activation_60_53), .reg_weight(reg_weight_60_53), .reg_partial_sum(reg_psum_60_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_54( .activation_in(reg_activation_60_53), .weight_in(reg_weight_59_54), .partial_sum_in(reg_psum_59_54), .reg_activation(reg_activation_60_54), .reg_weight(reg_weight_60_54), .reg_partial_sum(reg_psum_60_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_55( .activation_in(reg_activation_60_54), .weight_in(reg_weight_59_55), .partial_sum_in(reg_psum_59_55), .reg_activation(reg_activation_60_55), .reg_weight(reg_weight_60_55), .reg_partial_sum(reg_psum_60_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_56( .activation_in(reg_activation_60_55), .weight_in(reg_weight_59_56), .partial_sum_in(reg_psum_59_56), .reg_activation(reg_activation_60_56), .reg_weight(reg_weight_60_56), .reg_partial_sum(reg_psum_60_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_57( .activation_in(reg_activation_60_56), .weight_in(reg_weight_59_57), .partial_sum_in(reg_psum_59_57), .reg_activation(reg_activation_60_57), .reg_weight(reg_weight_60_57), .reg_partial_sum(reg_psum_60_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_58( .activation_in(reg_activation_60_57), .weight_in(reg_weight_59_58), .partial_sum_in(reg_psum_59_58), .reg_activation(reg_activation_60_58), .reg_weight(reg_weight_60_58), .reg_partial_sum(reg_psum_60_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_59( .activation_in(reg_activation_60_58), .weight_in(reg_weight_59_59), .partial_sum_in(reg_psum_59_59), .reg_activation(reg_activation_60_59), .reg_weight(reg_weight_60_59), .reg_partial_sum(reg_psum_60_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_60( .activation_in(reg_activation_60_59), .weight_in(reg_weight_59_60), .partial_sum_in(reg_psum_59_60), .reg_activation(reg_activation_60_60), .reg_weight(reg_weight_60_60), .reg_partial_sum(reg_psum_60_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_61( .activation_in(reg_activation_60_60), .weight_in(reg_weight_59_61), .partial_sum_in(reg_psum_59_61), .reg_activation(reg_activation_60_61), .reg_weight(reg_weight_60_61), .reg_partial_sum(reg_psum_60_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_62( .activation_in(reg_activation_60_61), .weight_in(reg_weight_59_62), .partial_sum_in(reg_psum_59_62), .reg_activation(reg_activation_60_62), .reg_weight(reg_weight_60_62), .reg_partial_sum(reg_psum_60_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U60_63( .activation_in(reg_activation_60_62), .weight_in(reg_weight_59_63), .partial_sum_in(reg_psum_59_63), .reg_weight(reg_weight_60_63), .reg_partial_sum(reg_psum_60_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_0( .activation_in(in_activation_61), .weight_in(reg_weight_60_0), .partial_sum_in(reg_psum_60_0), .reg_activation(reg_activation_61_0), .reg_weight(reg_weight_61_0), .reg_partial_sum(reg_psum_61_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_1( .activation_in(reg_activation_61_0), .weight_in(reg_weight_60_1), .partial_sum_in(reg_psum_60_1), .reg_activation(reg_activation_61_1), .reg_weight(reg_weight_61_1), .reg_partial_sum(reg_psum_61_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_2( .activation_in(reg_activation_61_1), .weight_in(reg_weight_60_2), .partial_sum_in(reg_psum_60_2), .reg_activation(reg_activation_61_2), .reg_weight(reg_weight_61_2), .reg_partial_sum(reg_psum_61_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_3( .activation_in(reg_activation_61_2), .weight_in(reg_weight_60_3), .partial_sum_in(reg_psum_60_3), .reg_activation(reg_activation_61_3), .reg_weight(reg_weight_61_3), .reg_partial_sum(reg_psum_61_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_4( .activation_in(reg_activation_61_3), .weight_in(reg_weight_60_4), .partial_sum_in(reg_psum_60_4), .reg_activation(reg_activation_61_4), .reg_weight(reg_weight_61_4), .reg_partial_sum(reg_psum_61_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_5( .activation_in(reg_activation_61_4), .weight_in(reg_weight_60_5), .partial_sum_in(reg_psum_60_5), .reg_activation(reg_activation_61_5), .reg_weight(reg_weight_61_5), .reg_partial_sum(reg_psum_61_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_6( .activation_in(reg_activation_61_5), .weight_in(reg_weight_60_6), .partial_sum_in(reg_psum_60_6), .reg_activation(reg_activation_61_6), .reg_weight(reg_weight_61_6), .reg_partial_sum(reg_psum_61_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_7( .activation_in(reg_activation_61_6), .weight_in(reg_weight_60_7), .partial_sum_in(reg_psum_60_7), .reg_activation(reg_activation_61_7), .reg_weight(reg_weight_61_7), .reg_partial_sum(reg_psum_61_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_8( .activation_in(reg_activation_61_7), .weight_in(reg_weight_60_8), .partial_sum_in(reg_psum_60_8), .reg_activation(reg_activation_61_8), .reg_weight(reg_weight_61_8), .reg_partial_sum(reg_psum_61_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_9( .activation_in(reg_activation_61_8), .weight_in(reg_weight_60_9), .partial_sum_in(reg_psum_60_9), .reg_activation(reg_activation_61_9), .reg_weight(reg_weight_61_9), .reg_partial_sum(reg_psum_61_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_10( .activation_in(reg_activation_61_9), .weight_in(reg_weight_60_10), .partial_sum_in(reg_psum_60_10), .reg_activation(reg_activation_61_10), .reg_weight(reg_weight_61_10), .reg_partial_sum(reg_psum_61_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_11( .activation_in(reg_activation_61_10), .weight_in(reg_weight_60_11), .partial_sum_in(reg_psum_60_11), .reg_activation(reg_activation_61_11), .reg_weight(reg_weight_61_11), .reg_partial_sum(reg_psum_61_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_12( .activation_in(reg_activation_61_11), .weight_in(reg_weight_60_12), .partial_sum_in(reg_psum_60_12), .reg_activation(reg_activation_61_12), .reg_weight(reg_weight_61_12), .reg_partial_sum(reg_psum_61_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_13( .activation_in(reg_activation_61_12), .weight_in(reg_weight_60_13), .partial_sum_in(reg_psum_60_13), .reg_activation(reg_activation_61_13), .reg_weight(reg_weight_61_13), .reg_partial_sum(reg_psum_61_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_14( .activation_in(reg_activation_61_13), .weight_in(reg_weight_60_14), .partial_sum_in(reg_psum_60_14), .reg_activation(reg_activation_61_14), .reg_weight(reg_weight_61_14), .reg_partial_sum(reg_psum_61_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_15( .activation_in(reg_activation_61_14), .weight_in(reg_weight_60_15), .partial_sum_in(reg_psum_60_15), .reg_activation(reg_activation_61_15), .reg_weight(reg_weight_61_15), .reg_partial_sum(reg_psum_61_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_16( .activation_in(reg_activation_61_15), .weight_in(reg_weight_60_16), .partial_sum_in(reg_psum_60_16), .reg_activation(reg_activation_61_16), .reg_weight(reg_weight_61_16), .reg_partial_sum(reg_psum_61_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_17( .activation_in(reg_activation_61_16), .weight_in(reg_weight_60_17), .partial_sum_in(reg_psum_60_17), .reg_activation(reg_activation_61_17), .reg_weight(reg_weight_61_17), .reg_partial_sum(reg_psum_61_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_18( .activation_in(reg_activation_61_17), .weight_in(reg_weight_60_18), .partial_sum_in(reg_psum_60_18), .reg_activation(reg_activation_61_18), .reg_weight(reg_weight_61_18), .reg_partial_sum(reg_psum_61_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_19( .activation_in(reg_activation_61_18), .weight_in(reg_weight_60_19), .partial_sum_in(reg_psum_60_19), .reg_activation(reg_activation_61_19), .reg_weight(reg_weight_61_19), .reg_partial_sum(reg_psum_61_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_20( .activation_in(reg_activation_61_19), .weight_in(reg_weight_60_20), .partial_sum_in(reg_psum_60_20), .reg_activation(reg_activation_61_20), .reg_weight(reg_weight_61_20), .reg_partial_sum(reg_psum_61_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_21( .activation_in(reg_activation_61_20), .weight_in(reg_weight_60_21), .partial_sum_in(reg_psum_60_21), .reg_activation(reg_activation_61_21), .reg_weight(reg_weight_61_21), .reg_partial_sum(reg_psum_61_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_22( .activation_in(reg_activation_61_21), .weight_in(reg_weight_60_22), .partial_sum_in(reg_psum_60_22), .reg_activation(reg_activation_61_22), .reg_weight(reg_weight_61_22), .reg_partial_sum(reg_psum_61_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_23( .activation_in(reg_activation_61_22), .weight_in(reg_weight_60_23), .partial_sum_in(reg_psum_60_23), .reg_activation(reg_activation_61_23), .reg_weight(reg_weight_61_23), .reg_partial_sum(reg_psum_61_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_24( .activation_in(reg_activation_61_23), .weight_in(reg_weight_60_24), .partial_sum_in(reg_psum_60_24), .reg_activation(reg_activation_61_24), .reg_weight(reg_weight_61_24), .reg_partial_sum(reg_psum_61_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_25( .activation_in(reg_activation_61_24), .weight_in(reg_weight_60_25), .partial_sum_in(reg_psum_60_25), .reg_activation(reg_activation_61_25), .reg_weight(reg_weight_61_25), .reg_partial_sum(reg_psum_61_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_26( .activation_in(reg_activation_61_25), .weight_in(reg_weight_60_26), .partial_sum_in(reg_psum_60_26), .reg_activation(reg_activation_61_26), .reg_weight(reg_weight_61_26), .reg_partial_sum(reg_psum_61_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_27( .activation_in(reg_activation_61_26), .weight_in(reg_weight_60_27), .partial_sum_in(reg_psum_60_27), .reg_activation(reg_activation_61_27), .reg_weight(reg_weight_61_27), .reg_partial_sum(reg_psum_61_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_28( .activation_in(reg_activation_61_27), .weight_in(reg_weight_60_28), .partial_sum_in(reg_psum_60_28), .reg_activation(reg_activation_61_28), .reg_weight(reg_weight_61_28), .reg_partial_sum(reg_psum_61_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_29( .activation_in(reg_activation_61_28), .weight_in(reg_weight_60_29), .partial_sum_in(reg_psum_60_29), .reg_activation(reg_activation_61_29), .reg_weight(reg_weight_61_29), .reg_partial_sum(reg_psum_61_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_30( .activation_in(reg_activation_61_29), .weight_in(reg_weight_60_30), .partial_sum_in(reg_psum_60_30), .reg_activation(reg_activation_61_30), .reg_weight(reg_weight_61_30), .reg_partial_sum(reg_psum_61_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_31( .activation_in(reg_activation_61_30), .weight_in(reg_weight_60_31), .partial_sum_in(reg_psum_60_31), .reg_activation(reg_activation_61_31), .reg_weight(reg_weight_61_31), .reg_partial_sum(reg_psum_61_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_32( .activation_in(reg_activation_61_31), .weight_in(reg_weight_60_32), .partial_sum_in(reg_psum_60_32), .reg_activation(reg_activation_61_32), .reg_weight(reg_weight_61_32), .reg_partial_sum(reg_psum_61_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_33( .activation_in(reg_activation_61_32), .weight_in(reg_weight_60_33), .partial_sum_in(reg_psum_60_33), .reg_activation(reg_activation_61_33), .reg_weight(reg_weight_61_33), .reg_partial_sum(reg_psum_61_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_34( .activation_in(reg_activation_61_33), .weight_in(reg_weight_60_34), .partial_sum_in(reg_psum_60_34), .reg_activation(reg_activation_61_34), .reg_weight(reg_weight_61_34), .reg_partial_sum(reg_psum_61_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_35( .activation_in(reg_activation_61_34), .weight_in(reg_weight_60_35), .partial_sum_in(reg_psum_60_35), .reg_activation(reg_activation_61_35), .reg_weight(reg_weight_61_35), .reg_partial_sum(reg_psum_61_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_36( .activation_in(reg_activation_61_35), .weight_in(reg_weight_60_36), .partial_sum_in(reg_psum_60_36), .reg_activation(reg_activation_61_36), .reg_weight(reg_weight_61_36), .reg_partial_sum(reg_psum_61_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_37( .activation_in(reg_activation_61_36), .weight_in(reg_weight_60_37), .partial_sum_in(reg_psum_60_37), .reg_activation(reg_activation_61_37), .reg_weight(reg_weight_61_37), .reg_partial_sum(reg_psum_61_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_38( .activation_in(reg_activation_61_37), .weight_in(reg_weight_60_38), .partial_sum_in(reg_psum_60_38), .reg_activation(reg_activation_61_38), .reg_weight(reg_weight_61_38), .reg_partial_sum(reg_psum_61_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_39( .activation_in(reg_activation_61_38), .weight_in(reg_weight_60_39), .partial_sum_in(reg_psum_60_39), .reg_activation(reg_activation_61_39), .reg_weight(reg_weight_61_39), .reg_partial_sum(reg_psum_61_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_40( .activation_in(reg_activation_61_39), .weight_in(reg_weight_60_40), .partial_sum_in(reg_psum_60_40), .reg_activation(reg_activation_61_40), .reg_weight(reg_weight_61_40), .reg_partial_sum(reg_psum_61_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_41( .activation_in(reg_activation_61_40), .weight_in(reg_weight_60_41), .partial_sum_in(reg_psum_60_41), .reg_activation(reg_activation_61_41), .reg_weight(reg_weight_61_41), .reg_partial_sum(reg_psum_61_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_42( .activation_in(reg_activation_61_41), .weight_in(reg_weight_60_42), .partial_sum_in(reg_psum_60_42), .reg_activation(reg_activation_61_42), .reg_weight(reg_weight_61_42), .reg_partial_sum(reg_psum_61_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_43( .activation_in(reg_activation_61_42), .weight_in(reg_weight_60_43), .partial_sum_in(reg_psum_60_43), .reg_activation(reg_activation_61_43), .reg_weight(reg_weight_61_43), .reg_partial_sum(reg_psum_61_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_44( .activation_in(reg_activation_61_43), .weight_in(reg_weight_60_44), .partial_sum_in(reg_psum_60_44), .reg_activation(reg_activation_61_44), .reg_weight(reg_weight_61_44), .reg_partial_sum(reg_psum_61_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_45( .activation_in(reg_activation_61_44), .weight_in(reg_weight_60_45), .partial_sum_in(reg_psum_60_45), .reg_activation(reg_activation_61_45), .reg_weight(reg_weight_61_45), .reg_partial_sum(reg_psum_61_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_46( .activation_in(reg_activation_61_45), .weight_in(reg_weight_60_46), .partial_sum_in(reg_psum_60_46), .reg_activation(reg_activation_61_46), .reg_weight(reg_weight_61_46), .reg_partial_sum(reg_psum_61_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_47( .activation_in(reg_activation_61_46), .weight_in(reg_weight_60_47), .partial_sum_in(reg_psum_60_47), .reg_activation(reg_activation_61_47), .reg_weight(reg_weight_61_47), .reg_partial_sum(reg_psum_61_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_48( .activation_in(reg_activation_61_47), .weight_in(reg_weight_60_48), .partial_sum_in(reg_psum_60_48), .reg_activation(reg_activation_61_48), .reg_weight(reg_weight_61_48), .reg_partial_sum(reg_psum_61_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_49( .activation_in(reg_activation_61_48), .weight_in(reg_weight_60_49), .partial_sum_in(reg_psum_60_49), .reg_activation(reg_activation_61_49), .reg_weight(reg_weight_61_49), .reg_partial_sum(reg_psum_61_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_50( .activation_in(reg_activation_61_49), .weight_in(reg_weight_60_50), .partial_sum_in(reg_psum_60_50), .reg_activation(reg_activation_61_50), .reg_weight(reg_weight_61_50), .reg_partial_sum(reg_psum_61_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_51( .activation_in(reg_activation_61_50), .weight_in(reg_weight_60_51), .partial_sum_in(reg_psum_60_51), .reg_activation(reg_activation_61_51), .reg_weight(reg_weight_61_51), .reg_partial_sum(reg_psum_61_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_52( .activation_in(reg_activation_61_51), .weight_in(reg_weight_60_52), .partial_sum_in(reg_psum_60_52), .reg_activation(reg_activation_61_52), .reg_weight(reg_weight_61_52), .reg_partial_sum(reg_psum_61_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_53( .activation_in(reg_activation_61_52), .weight_in(reg_weight_60_53), .partial_sum_in(reg_psum_60_53), .reg_activation(reg_activation_61_53), .reg_weight(reg_weight_61_53), .reg_partial_sum(reg_psum_61_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_54( .activation_in(reg_activation_61_53), .weight_in(reg_weight_60_54), .partial_sum_in(reg_psum_60_54), .reg_activation(reg_activation_61_54), .reg_weight(reg_weight_61_54), .reg_partial_sum(reg_psum_61_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_55( .activation_in(reg_activation_61_54), .weight_in(reg_weight_60_55), .partial_sum_in(reg_psum_60_55), .reg_activation(reg_activation_61_55), .reg_weight(reg_weight_61_55), .reg_partial_sum(reg_psum_61_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_56( .activation_in(reg_activation_61_55), .weight_in(reg_weight_60_56), .partial_sum_in(reg_psum_60_56), .reg_activation(reg_activation_61_56), .reg_weight(reg_weight_61_56), .reg_partial_sum(reg_psum_61_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_57( .activation_in(reg_activation_61_56), .weight_in(reg_weight_60_57), .partial_sum_in(reg_psum_60_57), .reg_activation(reg_activation_61_57), .reg_weight(reg_weight_61_57), .reg_partial_sum(reg_psum_61_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_58( .activation_in(reg_activation_61_57), .weight_in(reg_weight_60_58), .partial_sum_in(reg_psum_60_58), .reg_activation(reg_activation_61_58), .reg_weight(reg_weight_61_58), .reg_partial_sum(reg_psum_61_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_59( .activation_in(reg_activation_61_58), .weight_in(reg_weight_60_59), .partial_sum_in(reg_psum_60_59), .reg_activation(reg_activation_61_59), .reg_weight(reg_weight_61_59), .reg_partial_sum(reg_psum_61_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_60( .activation_in(reg_activation_61_59), .weight_in(reg_weight_60_60), .partial_sum_in(reg_psum_60_60), .reg_activation(reg_activation_61_60), .reg_weight(reg_weight_61_60), .reg_partial_sum(reg_psum_61_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_61( .activation_in(reg_activation_61_60), .weight_in(reg_weight_60_61), .partial_sum_in(reg_psum_60_61), .reg_activation(reg_activation_61_61), .reg_weight(reg_weight_61_61), .reg_partial_sum(reg_psum_61_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_62( .activation_in(reg_activation_61_61), .weight_in(reg_weight_60_62), .partial_sum_in(reg_psum_60_62), .reg_activation(reg_activation_61_62), .reg_weight(reg_weight_61_62), .reg_partial_sum(reg_psum_61_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U61_63( .activation_in(reg_activation_61_62), .weight_in(reg_weight_60_63), .partial_sum_in(reg_psum_60_63), .reg_weight(reg_weight_61_63), .reg_partial_sum(reg_psum_61_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_0( .activation_in(in_activation_62), .weight_in(reg_weight_61_0), .partial_sum_in(reg_psum_61_0), .reg_activation(reg_activation_62_0), .reg_weight(reg_weight_62_0), .reg_partial_sum(reg_psum_62_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_1( .activation_in(reg_activation_62_0), .weight_in(reg_weight_61_1), .partial_sum_in(reg_psum_61_1), .reg_activation(reg_activation_62_1), .reg_weight(reg_weight_62_1), .reg_partial_sum(reg_psum_62_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_2( .activation_in(reg_activation_62_1), .weight_in(reg_weight_61_2), .partial_sum_in(reg_psum_61_2), .reg_activation(reg_activation_62_2), .reg_weight(reg_weight_62_2), .reg_partial_sum(reg_psum_62_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_3( .activation_in(reg_activation_62_2), .weight_in(reg_weight_61_3), .partial_sum_in(reg_psum_61_3), .reg_activation(reg_activation_62_3), .reg_weight(reg_weight_62_3), .reg_partial_sum(reg_psum_62_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_4( .activation_in(reg_activation_62_3), .weight_in(reg_weight_61_4), .partial_sum_in(reg_psum_61_4), .reg_activation(reg_activation_62_4), .reg_weight(reg_weight_62_4), .reg_partial_sum(reg_psum_62_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_5( .activation_in(reg_activation_62_4), .weight_in(reg_weight_61_5), .partial_sum_in(reg_psum_61_5), .reg_activation(reg_activation_62_5), .reg_weight(reg_weight_62_5), .reg_partial_sum(reg_psum_62_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_6( .activation_in(reg_activation_62_5), .weight_in(reg_weight_61_6), .partial_sum_in(reg_psum_61_6), .reg_activation(reg_activation_62_6), .reg_weight(reg_weight_62_6), .reg_partial_sum(reg_psum_62_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_7( .activation_in(reg_activation_62_6), .weight_in(reg_weight_61_7), .partial_sum_in(reg_psum_61_7), .reg_activation(reg_activation_62_7), .reg_weight(reg_weight_62_7), .reg_partial_sum(reg_psum_62_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_8( .activation_in(reg_activation_62_7), .weight_in(reg_weight_61_8), .partial_sum_in(reg_psum_61_8), .reg_activation(reg_activation_62_8), .reg_weight(reg_weight_62_8), .reg_partial_sum(reg_psum_62_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_9( .activation_in(reg_activation_62_8), .weight_in(reg_weight_61_9), .partial_sum_in(reg_psum_61_9), .reg_activation(reg_activation_62_9), .reg_weight(reg_weight_62_9), .reg_partial_sum(reg_psum_62_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_10( .activation_in(reg_activation_62_9), .weight_in(reg_weight_61_10), .partial_sum_in(reg_psum_61_10), .reg_activation(reg_activation_62_10), .reg_weight(reg_weight_62_10), .reg_partial_sum(reg_psum_62_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_11( .activation_in(reg_activation_62_10), .weight_in(reg_weight_61_11), .partial_sum_in(reg_psum_61_11), .reg_activation(reg_activation_62_11), .reg_weight(reg_weight_62_11), .reg_partial_sum(reg_psum_62_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_12( .activation_in(reg_activation_62_11), .weight_in(reg_weight_61_12), .partial_sum_in(reg_psum_61_12), .reg_activation(reg_activation_62_12), .reg_weight(reg_weight_62_12), .reg_partial_sum(reg_psum_62_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_13( .activation_in(reg_activation_62_12), .weight_in(reg_weight_61_13), .partial_sum_in(reg_psum_61_13), .reg_activation(reg_activation_62_13), .reg_weight(reg_weight_62_13), .reg_partial_sum(reg_psum_62_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_14( .activation_in(reg_activation_62_13), .weight_in(reg_weight_61_14), .partial_sum_in(reg_psum_61_14), .reg_activation(reg_activation_62_14), .reg_weight(reg_weight_62_14), .reg_partial_sum(reg_psum_62_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_15( .activation_in(reg_activation_62_14), .weight_in(reg_weight_61_15), .partial_sum_in(reg_psum_61_15), .reg_activation(reg_activation_62_15), .reg_weight(reg_weight_62_15), .reg_partial_sum(reg_psum_62_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_16( .activation_in(reg_activation_62_15), .weight_in(reg_weight_61_16), .partial_sum_in(reg_psum_61_16), .reg_activation(reg_activation_62_16), .reg_weight(reg_weight_62_16), .reg_partial_sum(reg_psum_62_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_17( .activation_in(reg_activation_62_16), .weight_in(reg_weight_61_17), .partial_sum_in(reg_psum_61_17), .reg_activation(reg_activation_62_17), .reg_weight(reg_weight_62_17), .reg_partial_sum(reg_psum_62_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_18( .activation_in(reg_activation_62_17), .weight_in(reg_weight_61_18), .partial_sum_in(reg_psum_61_18), .reg_activation(reg_activation_62_18), .reg_weight(reg_weight_62_18), .reg_partial_sum(reg_psum_62_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_19( .activation_in(reg_activation_62_18), .weight_in(reg_weight_61_19), .partial_sum_in(reg_psum_61_19), .reg_activation(reg_activation_62_19), .reg_weight(reg_weight_62_19), .reg_partial_sum(reg_psum_62_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_20( .activation_in(reg_activation_62_19), .weight_in(reg_weight_61_20), .partial_sum_in(reg_psum_61_20), .reg_activation(reg_activation_62_20), .reg_weight(reg_weight_62_20), .reg_partial_sum(reg_psum_62_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_21( .activation_in(reg_activation_62_20), .weight_in(reg_weight_61_21), .partial_sum_in(reg_psum_61_21), .reg_activation(reg_activation_62_21), .reg_weight(reg_weight_62_21), .reg_partial_sum(reg_psum_62_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_22( .activation_in(reg_activation_62_21), .weight_in(reg_weight_61_22), .partial_sum_in(reg_psum_61_22), .reg_activation(reg_activation_62_22), .reg_weight(reg_weight_62_22), .reg_partial_sum(reg_psum_62_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_23( .activation_in(reg_activation_62_22), .weight_in(reg_weight_61_23), .partial_sum_in(reg_psum_61_23), .reg_activation(reg_activation_62_23), .reg_weight(reg_weight_62_23), .reg_partial_sum(reg_psum_62_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_24( .activation_in(reg_activation_62_23), .weight_in(reg_weight_61_24), .partial_sum_in(reg_psum_61_24), .reg_activation(reg_activation_62_24), .reg_weight(reg_weight_62_24), .reg_partial_sum(reg_psum_62_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_25( .activation_in(reg_activation_62_24), .weight_in(reg_weight_61_25), .partial_sum_in(reg_psum_61_25), .reg_activation(reg_activation_62_25), .reg_weight(reg_weight_62_25), .reg_partial_sum(reg_psum_62_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_26( .activation_in(reg_activation_62_25), .weight_in(reg_weight_61_26), .partial_sum_in(reg_psum_61_26), .reg_activation(reg_activation_62_26), .reg_weight(reg_weight_62_26), .reg_partial_sum(reg_psum_62_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_27( .activation_in(reg_activation_62_26), .weight_in(reg_weight_61_27), .partial_sum_in(reg_psum_61_27), .reg_activation(reg_activation_62_27), .reg_weight(reg_weight_62_27), .reg_partial_sum(reg_psum_62_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_28( .activation_in(reg_activation_62_27), .weight_in(reg_weight_61_28), .partial_sum_in(reg_psum_61_28), .reg_activation(reg_activation_62_28), .reg_weight(reg_weight_62_28), .reg_partial_sum(reg_psum_62_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_29( .activation_in(reg_activation_62_28), .weight_in(reg_weight_61_29), .partial_sum_in(reg_psum_61_29), .reg_activation(reg_activation_62_29), .reg_weight(reg_weight_62_29), .reg_partial_sum(reg_psum_62_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_30( .activation_in(reg_activation_62_29), .weight_in(reg_weight_61_30), .partial_sum_in(reg_psum_61_30), .reg_activation(reg_activation_62_30), .reg_weight(reg_weight_62_30), .reg_partial_sum(reg_psum_62_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_31( .activation_in(reg_activation_62_30), .weight_in(reg_weight_61_31), .partial_sum_in(reg_psum_61_31), .reg_activation(reg_activation_62_31), .reg_weight(reg_weight_62_31), .reg_partial_sum(reg_psum_62_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_32( .activation_in(reg_activation_62_31), .weight_in(reg_weight_61_32), .partial_sum_in(reg_psum_61_32), .reg_activation(reg_activation_62_32), .reg_weight(reg_weight_62_32), .reg_partial_sum(reg_psum_62_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_33( .activation_in(reg_activation_62_32), .weight_in(reg_weight_61_33), .partial_sum_in(reg_psum_61_33), .reg_activation(reg_activation_62_33), .reg_weight(reg_weight_62_33), .reg_partial_sum(reg_psum_62_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_34( .activation_in(reg_activation_62_33), .weight_in(reg_weight_61_34), .partial_sum_in(reg_psum_61_34), .reg_activation(reg_activation_62_34), .reg_weight(reg_weight_62_34), .reg_partial_sum(reg_psum_62_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_35( .activation_in(reg_activation_62_34), .weight_in(reg_weight_61_35), .partial_sum_in(reg_psum_61_35), .reg_activation(reg_activation_62_35), .reg_weight(reg_weight_62_35), .reg_partial_sum(reg_psum_62_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_36( .activation_in(reg_activation_62_35), .weight_in(reg_weight_61_36), .partial_sum_in(reg_psum_61_36), .reg_activation(reg_activation_62_36), .reg_weight(reg_weight_62_36), .reg_partial_sum(reg_psum_62_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_37( .activation_in(reg_activation_62_36), .weight_in(reg_weight_61_37), .partial_sum_in(reg_psum_61_37), .reg_activation(reg_activation_62_37), .reg_weight(reg_weight_62_37), .reg_partial_sum(reg_psum_62_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_38( .activation_in(reg_activation_62_37), .weight_in(reg_weight_61_38), .partial_sum_in(reg_psum_61_38), .reg_activation(reg_activation_62_38), .reg_weight(reg_weight_62_38), .reg_partial_sum(reg_psum_62_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_39( .activation_in(reg_activation_62_38), .weight_in(reg_weight_61_39), .partial_sum_in(reg_psum_61_39), .reg_activation(reg_activation_62_39), .reg_weight(reg_weight_62_39), .reg_partial_sum(reg_psum_62_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_40( .activation_in(reg_activation_62_39), .weight_in(reg_weight_61_40), .partial_sum_in(reg_psum_61_40), .reg_activation(reg_activation_62_40), .reg_weight(reg_weight_62_40), .reg_partial_sum(reg_psum_62_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_41( .activation_in(reg_activation_62_40), .weight_in(reg_weight_61_41), .partial_sum_in(reg_psum_61_41), .reg_activation(reg_activation_62_41), .reg_weight(reg_weight_62_41), .reg_partial_sum(reg_psum_62_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_42( .activation_in(reg_activation_62_41), .weight_in(reg_weight_61_42), .partial_sum_in(reg_psum_61_42), .reg_activation(reg_activation_62_42), .reg_weight(reg_weight_62_42), .reg_partial_sum(reg_psum_62_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_43( .activation_in(reg_activation_62_42), .weight_in(reg_weight_61_43), .partial_sum_in(reg_psum_61_43), .reg_activation(reg_activation_62_43), .reg_weight(reg_weight_62_43), .reg_partial_sum(reg_psum_62_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_44( .activation_in(reg_activation_62_43), .weight_in(reg_weight_61_44), .partial_sum_in(reg_psum_61_44), .reg_activation(reg_activation_62_44), .reg_weight(reg_weight_62_44), .reg_partial_sum(reg_psum_62_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_45( .activation_in(reg_activation_62_44), .weight_in(reg_weight_61_45), .partial_sum_in(reg_psum_61_45), .reg_activation(reg_activation_62_45), .reg_weight(reg_weight_62_45), .reg_partial_sum(reg_psum_62_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_46( .activation_in(reg_activation_62_45), .weight_in(reg_weight_61_46), .partial_sum_in(reg_psum_61_46), .reg_activation(reg_activation_62_46), .reg_weight(reg_weight_62_46), .reg_partial_sum(reg_psum_62_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_47( .activation_in(reg_activation_62_46), .weight_in(reg_weight_61_47), .partial_sum_in(reg_psum_61_47), .reg_activation(reg_activation_62_47), .reg_weight(reg_weight_62_47), .reg_partial_sum(reg_psum_62_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_48( .activation_in(reg_activation_62_47), .weight_in(reg_weight_61_48), .partial_sum_in(reg_psum_61_48), .reg_activation(reg_activation_62_48), .reg_weight(reg_weight_62_48), .reg_partial_sum(reg_psum_62_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_49( .activation_in(reg_activation_62_48), .weight_in(reg_weight_61_49), .partial_sum_in(reg_psum_61_49), .reg_activation(reg_activation_62_49), .reg_weight(reg_weight_62_49), .reg_partial_sum(reg_psum_62_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_50( .activation_in(reg_activation_62_49), .weight_in(reg_weight_61_50), .partial_sum_in(reg_psum_61_50), .reg_activation(reg_activation_62_50), .reg_weight(reg_weight_62_50), .reg_partial_sum(reg_psum_62_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_51( .activation_in(reg_activation_62_50), .weight_in(reg_weight_61_51), .partial_sum_in(reg_psum_61_51), .reg_activation(reg_activation_62_51), .reg_weight(reg_weight_62_51), .reg_partial_sum(reg_psum_62_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_52( .activation_in(reg_activation_62_51), .weight_in(reg_weight_61_52), .partial_sum_in(reg_psum_61_52), .reg_activation(reg_activation_62_52), .reg_weight(reg_weight_62_52), .reg_partial_sum(reg_psum_62_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_53( .activation_in(reg_activation_62_52), .weight_in(reg_weight_61_53), .partial_sum_in(reg_psum_61_53), .reg_activation(reg_activation_62_53), .reg_weight(reg_weight_62_53), .reg_partial_sum(reg_psum_62_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_54( .activation_in(reg_activation_62_53), .weight_in(reg_weight_61_54), .partial_sum_in(reg_psum_61_54), .reg_activation(reg_activation_62_54), .reg_weight(reg_weight_62_54), .reg_partial_sum(reg_psum_62_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_55( .activation_in(reg_activation_62_54), .weight_in(reg_weight_61_55), .partial_sum_in(reg_psum_61_55), .reg_activation(reg_activation_62_55), .reg_weight(reg_weight_62_55), .reg_partial_sum(reg_psum_62_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_56( .activation_in(reg_activation_62_55), .weight_in(reg_weight_61_56), .partial_sum_in(reg_psum_61_56), .reg_activation(reg_activation_62_56), .reg_weight(reg_weight_62_56), .reg_partial_sum(reg_psum_62_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_57( .activation_in(reg_activation_62_56), .weight_in(reg_weight_61_57), .partial_sum_in(reg_psum_61_57), .reg_activation(reg_activation_62_57), .reg_weight(reg_weight_62_57), .reg_partial_sum(reg_psum_62_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_58( .activation_in(reg_activation_62_57), .weight_in(reg_weight_61_58), .partial_sum_in(reg_psum_61_58), .reg_activation(reg_activation_62_58), .reg_weight(reg_weight_62_58), .reg_partial_sum(reg_psum_62_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_59( .activation_in(reg_activation_62_58), .weight_in(reg_weight_61_59), .partial_sum_in(reg_psum_61_59), .reg_activation(reg_activation_62_59), .reg_weight(reg_weight_62_59), .reg_partial_sum(reg_psum_62_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_60( .activation_in(reg_activation_62_59), .weight_in(reg_weight_61_60), .partial_sum_in(reg_psum_61_60), .reg_activation(reg_activation_62_60), .reg_weight(reg_weight_62_60), .reg_partial_sum(reg_psum_62_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_61( .activation_in(reg_activation_62_60), .weight_in(reg_weight_61_61), .partial_sum_in(reg_psum_61_61), .reg_activation(reg_activation_62_61), .reg_weight(reg_weight_62_61), .reg_partial_sum(reg_psum_62_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_62( .activation_in(reg_activation_62_61), .weight_in(reg_weight_61_62), .partial_sum_in(reg_psum_61_62), .reg_activation(reg_activation_62_62), .reg_weight(reg_weight_62_62), .reg_partial_sum(reg_psum_62_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U62_63( .activation_in(reg_activation_62_62), .weight_in(reg_weight_61_63), .partial_sum_in(reg_psum_61_63), .reg_weight(reg_weight_62_63), .reg_partial_sum(reg_psum_62_63), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_0( .activation_in(in_activation_63), .weight_in(reg_weight_62_0), .partial_sum_in(reg_psum_62_0), .reg_activation(reg_activation_63_0), .reg_partial_sum(reg_psum_63_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_1( .activation_in(reg_activation_63_0), .weight_in(reg_weight_62_1), .partial_sum_in(reg_psum_62_1), .reg_activation(reg_activation_63_1), .reg_partial_sum(reg_psum_63_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_2( .activation_in(reg_activation_63_1), .weight_in(reg_weight_62_2), .partial_sum_in(reg_psum_62_2), .reg_activation(reg_activation_63_2), .reg_partial_sum(reg_psum_63_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_3( .activation_in(reg_activation_63_2), .weight_in(reg_weight_62_3), .partial_sum_in(reg_psum_62_3), .reg_activation(reg_activation_63_3), .reg_partial_sum(reg_psum_63_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_4( .activation_in(reg_activation_63_3), .weight_in(reg_weight_62_4), .partial_sum_in(reg_psum_62_4), .reg_activation(reg_activation_63_4), .reg_partial_sum(reg_psum_63_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_5( .activation_in(reg_activation_63_4), .weight_in(reg_weight_62_5), .partial_sum_in(reg_psum_62_5), .reg_activation(reg_activation_63_5), .reg_partial_sum(reg_psum_63_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_6( .activation_in(reg_activation_63_5), .weight_in(reg_weight_62_6), .partial_sum_in(reg_psum_62_6), .reg_activation(reg_activation_63_6), .reg_partial_sum(reg_psum_63_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_7( .activation_in(reg_activation_63_6), .weight_in(reg_weight_62_7), .partial_sum_in(reg_psum_62_7), .reg_activation(reg_activation_63_7), .reg_partial_sum(reg_psum_63_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_8( .activation_in(reg_activation_63_7), .weight_in(reg_weight_62_8), .partial_sum_in(reg_psum_62_8), .reg_activation(reg_activation_63_8), .reg_partial_sum(reg_psum_63_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_9( .activation_in(reg_activation_63_8), .weight_in(reg_weight_62_9), .partial_sum_in(reg_psum_62_9), .reg_activation(reg_activation_63_9), .reg_partial_sum(reg_psum_63_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_10( .activation_in(reg_activation_63_9), .weight_in(reg_weight_62_10), .partial_sum_in(reg_psum_62_10), .reg_activation(reg_activation_63_10), .reg_partial_sum(reg_psum_63_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_11( .activation_in(reg_activation_63_10), .weight_in(reg_weight_62_11), .partial_sum_in(reg_psum_62_11), .reg_activation(reg_activation_63_11), .reg_partial_sum(reg_psum_63_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_12( .activation_in(reg_activation_63_11), .weight_in(reg_weight_62_12), .partial_sum_in(reg_psum_62_12), .reg_activation(reg_activation_63_12), .reg_partial_sum(reg_psum_63_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_13( .activation_in(reg_activation_63_12), .weight_in(reg_weight_62_13), .partial_sum_in(reg_psum_62_13), .reg_activation(reg_activation_63_13), .reg_partial_sum(reg_psum_63_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_14( .activation_in(reg_activation_63_13), .weight_in(reg_weight_62_14), .partial_sum_in(reg_psum_62_14), .reg_activation(reg_activation_63_14), .reg_partial_sum(reg_psum_63_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_15( .activation_in(reg_activation_63_14), .weight_in(reg_weight_62_15), .partial_sum_in(reg_psum_62_15), .reg_activation(reg_activation_63_15), .reg_partial_sum(reg_psum_63_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_16( .activation_in(reg_activation_63_15), .weight_in(reg_weight_62_16), .partial_sum_in(reg_psum_62_16), .reg_activation(reg_activation_63_16), .reg_partial_sum(reg_psum_63_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_17( .activation_in(reg_activation_63_16), .weight_in(reg_weight_62_17), .partial_sum_in(reg_psum_62_17), .reg_activation(reg_activation_63_17), .reg_partial_sum(reg_psum_63_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_18( .activation_in(reg_activation_63_17), .weight_in(reg_weight_62_18), .partial_sum_in(reg_psum_62_18), .reg_activation(reg_activation_63_18), .reg_partial_sum(reg_psum_63_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_19( .activation_in(reg_activation_63_18), .weight_in(reg_weight_62_19), .partial_sum_in(reg_psum_62_19), .reg_activation(reg_activation_63_19), .reg_partial_sum(reg_psum_63_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_20( .activation_in(reg_activation_63_19), .weight_in(reg_weight_62_20), .partial_sum_in(reg_psum_62_20), .reg_activation(reg_activation_63_20), .reg_partial_sum(reg_psum_63_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_21( .activation_in(reg_activation_63_20), .weight_in(reg_weight_62_21), .partial_sum_in(reg_psum_62_21), .reg_activation(reg_activation_63_21), .reg_partial_sum(reg_psum_63_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_22( .activation_in(reg_activation_63_21), .weight_in(reg_weight_62_22), .partial_sum_in(reg_psum_62_22), .reg_activation(reg_activation_63_22), .reg_partial_sum(reg_psum_63_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_23( .activation_in(reg_activation_63_22), .weight_in(reg_weight_62_23), .partial_sum_in(reg_psum_62_23), .reg_activation(reg_activation_63_23), .reg_partial_sum(reg_psum_63_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_24( .activation_in(reg_activation_63_23), .weight_in(reg_weight_62_24), .partial_sum_in(reg_psum_62_24), .reg_activation(reg_activation_63_24), .reg_partial_sum(reg_psum_63_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_25( .activation_in(reg_activation_63_24), .weight_in(reg_weight_62_25), .partial_sum_in(reg_psum_62_25), .reg_activation(reg_activation_63_25), .reg_partial_sum(reg_psum_63_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_26( .activation_in(reg_activation_63_25), .weight_in(reg_weight_62_26), .partial_sum_in(reg_psum_62_26), .reg_activation(reg_activation_63_26), .reg_partial_sum(reg_psum_63_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_27( .activation_in(reg_activation_63_26), .weight_in(reg_weight_62_27), .partial_sum_in(reg_psum_62_27), .reg_activation(reg_activation_63_27), .reg_partial_sum(reg_psum_63_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_28( .activation_in(reg_activation_63_27), .weight_in(reg_weight_62_28), .partial_sum_in(reg_psum_62_28), .reg_activation(reg_activation_63_28), .reg_partial_sum(reg_psum_63_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_29( .activation_in(reg_activation_63_28), .weight_in(reg_weight_62_29), .partial_sum_in(reg_psum_62_29), .reg_activation(reg_activation_63_29), .reg_partial_sum(reg_psum_63_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_30( .activation_in(reg_activation_63_29), .weight_in(reg_weight_62_30), .partial_sum_in(reg_psum_62_30), .reg_activation(reg_activation_63_30), .reg_partial_sum(reg_psum_63_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_31( .activation_in(reg_activation_63_30), .weight_in(reg_weight_62_31), .partial_sum_in(reg_psum_62_31), .reg_activation(reg_activation_63_31), .reg_partial_sum(reg_psum_63_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_32( .activation_in(reg_activation_63_31), .weight_in(reg_weight_62_32), .partial_sum_in(reg_psum_62_32), .reg_activation(reg_activation_63_32), .reg_partial_sum(reg_psum_63_32), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_33( .activation_in(reg_activation_63_32), .weight_in(reg_weight_62_33), .partial_sum_in(reg_psum_62_33), .reg_activation(reg_activation_63_33), .reg_partial_sum(reg_psum_63_33), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_34( .activation_in(reg_activation_63_33), .weight_in(reg_weight_62_34), .partial_sum_in(reg_psum_62_34), .reg_activation(reg_activation_63_34), .reg_partial_sum(reg_psum_63_34), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_35( .activation_in(reg_activation_63_34), .weight_in(reg_weight_62_35), .partial_sum_in(reg_psum_62_35), .reg_activation(reg_activation_63_35), .reg_partial_sum(reg_psum_63_35), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_36( .activation_in(reg_activation_63_35), .weight_in(reg_weight_62_36), .partial_sum_in(reg_psum_62_36), .reg_activation(reg_activation_63_36), .reg_partial_sum(reg_psum_63_36), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_37( .activation_in(reg_activation_63_36), .weight_in(reg_weight_62_37), .partial_sum_in(reg_psum_62_37), .reg_activation(reg_activation_63_37), .reg_partial_sum(reg_psum_63_37), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_38( .activation_in(reg_activation_63_37), .weight_in(reg_weight_62_38), .partial_sum_in(reg_psum_62_38), .reg_activation(reg_activation_63_38), .reg_partial_sum(reg_psum_63_38), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_39( .activation_in(reg_activation_63_38), .weight_in(reg_weight_62_39), .partial_sum_in(reg_psum_62_39), .reg_activation(reg_activation_63_39), .reg_partial_sum(reg_psum_63_39), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_40( .activation_in(reg_activation_63_39), .weight_in(reg_weight_62_40), .partial_sum_in(reg_psum_62_40), .reg_activation(reg_activation_63_40), .reg_partial_sum(reg_psum_63_40), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_41( .activation_in(reg_activation_63_40), .weight_in(reg_weight_62_41), .partial_sum_in(reg_psum_62_41), .reg_activation(reg_activation_63_41), .reg_partial_sum(reg_psum_63_41), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_42( .activation_in(reg_activation_63_41), .weight_in(reg_weight_62_42), .partial_sum_in(reg_psum_62_42), .reg_activation(reg_activation_63_42), .reg_partial_sum(reg_psum_63_42), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_43( .activation_in(reg_activation_63_42), .weight_in(reg_weight_62_43), .partial_sum_in(reg_psum_62_43), .reg_activation(reg_activation_63_43), .reg_partial_sum(reg_psum_63_43), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_44( .activation_in(reg_activation_63_43), .weight_in(reg_weight_62_44), .partial_sum_in(reg_psum_62_44), .reg_activation(reg_activation_63_44), .reg_partial_sum(reg_psum_63_44), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_45( .activation_in(reg_activation_63_44), .weight_in(reg_weight_62_45), .partial_sum_in(reg_psum_62_45), .reg_activation(reg_activation_63_45), .reg_partial_sum(reg_psum_63_45), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_46( .activation_in(reg_activation_63_45), .weight_in(reg_weight_62_46), .partial_sum_in(reg_psum_62_46), .reg_activation(reg_activation_63_46), .reg_partial_sum(reg_psum_63_46), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_47( .activation_in(reg_activation_63_46), .weight_in(reg_weight_62_47), .partial_sum_in(reg_psum_62_47), .reg_activation(reg_activation_63_47), .reg_partial_sum(reg_psum_63_47), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_48( .activation_in(reg_activation_63_47), .weight_in(reg_weight_62_48), .partial_sum_in(reg_psum_62_48), .reg_activation(reg_activation_63_48), .reg_partial_sum(reg_psum_63_48), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_49( .activation_in(reg_activation_63_48), .weight_in(reg_weight_62_49), .partial_sum_in(reg_psum_62_49), .reg_activation(reg_activation_63_49), .reg_partial_sum(reg_psum_63_49), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_50( .activation_in(reg_activation_63_49), .weight_in(reg_weight_62_50), .partial_sum_in(reg_psum_62_50), .reg_activation(reg_activation_63_50), .reg_partial_sum(reg_psum_63_50), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_51( .activation_in(reg_activation_63_50), .weight_in(reg_weight_62_51), .partial_sum_in(reg_psum_62_51), .reg_activation(reg_activation_63_51), .reg_partial_sum(reg_psum_63_51), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_52( .activation_in(reg_activation_63_51), .weight_in(reg_weight_62_52), .partial_sum_in(reg_psum_62_52), .reg_activation(reg_activation_63_52), .reg_partial_sum(reg_psum_63_52), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_53( .activation_in(reg_activation_63_52), .weight_in(reg_weight_62_53), .partial_sum_in(reg_psum_62_53), .reg_activation(reg_activation_63_53), .reg_partial_sum(reg_psum_63_53), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_54( .activation_in(reg_activation_63_53), .weight_in(reg_weight_62_54), .partial_sum_in(reg_psum_62_54), .reg_activation(reg_activation_63_54), .reg_partial_sum(reg_psum_63_54), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_55( .activation_in(reg_activation_63_54), .weight_in(reg_weight_62_55), .partial_sum_in(reg_psum_62_55), .reg_activation(reg_activation_63_55), .reg_partial_sum(reg_psum_63_55), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_56( .activation_in(reg_activation_63_55), .weight_in(reg_weight_62_56), .partial_sum_in(reg_psum_62_56), .reg_activation(reg_activation_63_56), .reg_partial_sum(reg_psum_63_56), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_57( .activation_in(reg_activation_63_56), .weight_in(reg_weight_62_57), .partial_sum_in(reg_psum_62_57), .reg_activation(reg_activation_63_57), .reg_partial_sum(reg_psum_63_57), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_58( .activation_in(reg_activation_63_57), .weight_in(reg_weight_62_58), .partial_sum_in(reg_psum_62_58), .reg_activation(reg_activation_63_58), .reg_partial_sum(reg_psum_63_58), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_59( .activation_in(reg_activation_63_58), .weight_in(reg_weight_62_59), .partial_sum_in(reg_psum_62_59), .reg_activation(reg_activation_63_59), .reg_partial_sum(reg_psum_63_59), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_60( .activation_in(reg_activation_63_59), .weight_in(reg_weight_62_60), .partial_sum_in(reg_psum_62_60), .reg_activation(reg_activation_63_60), .reg_partial_sum(reg_psum_63_60), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_61( .activation_in(reg_activation_63_60), .weight_in(reg_weight_62_61), .partial_sum_in(reg_psum_62_61), .reg_activation(reg_activation_63_61), .reg_partial_sum(reg_psum_63_61), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_62( .activation_in(reg_activation_63_61), .weight_in(reg_weight_62_62), .partial_sum_in(reg_psum_62_62), .reg_activation(reg_activation_63_62), .reg_partial_sum(reg_psum_63_62), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U63_63( .activation_in(reg_activation_63_62), .weight_in(reg_weight_62_63), .partial_sum_in(reg_psum_62_63), .reg_partial_sum(reg_psum_63_63), .clk(clk), .rst(rst), .weight_en(weight_en));
assign out_psum_0 = reg_psum_63_0;
assign out_psum_1 = reg_psum_63_1;
assign out_psum_2 = reg_psum_63_2;
assign out_psum_3 = reg_psum_63_3;
assign out_psum_4 = reg_psum_63_4;
assign out_psum_5 = reg_psum_63_5;
assign out_psum_6 = reg_psum_63_6;
assign out_psum_7 = reg_psum_63_7;
assign out_psum_8 = reg_psum_63_8;
assign out_psum_9 = reg_psum_63_9;
assign out_psum_10 = reg_psum_63_10;
assign out_psum_11 = reg_psum_63_11;
assign out_psum_12 = reg_psum_63_12;
assign out_psum_13 = reg_psum_63_13;
assign out_psum_14 = reg_psum_63_14;
assign out_psum_15 = reg_psum_63_15;
assign out_psum_16 = reg_psum_63_16;
assign out_psum_17 = reg_psum_63_17;
assign out_psum_18 = reg_psum_63_18;
assign out_psum_19 = reg_psum_63_19;
assign out_psum_20 = reg_psum_63_20;
assign out_psum_21 = reg_psum_63_21;
assign out_psum_22 = reg_psum_63_22;
assign out_psum_23 = reg_psum_63_23;
assign out_psum_24 = reg_psum_63_24;
assign out_psum_25 = reg_psum_63_25;
assign out_psum_26 = reg_psum_63_26;
assign out_psum_27 = reg_psum_63_27;
assign out_psum_28 = reg_psum_63_28;
assign out_psum_29 = reg_psum_63_29;
assign out_psum_30 = reg_psum_63_30;
assign out_psum_31 = reg_psum_63_31;
assign out_psum_32 = reg_psum_63_32;
assign out_psum_33 = reg_psum_63_33;
assign out_psum_34 = reg_psum_63_34;
assign out_psum_35 = reg_psum_63_35;
assign out_psum_36 = reg_psum_63_36;
assign out_psum_37 = reg_psum_63_37;
assign out_psum_38 = reg_psum_63_38;
assign out_psum_39 = reg_psum_63_39;
assign out_psum_40 = reg_psum_63_40;
assign out_psum_41 = reg_psum_63_41;
assign out_psum_42 = reg_psum_63_42;
assign out_psum_43 = reg_psum_63_43;
assign out_psum_44 = reg_psum_63_44;
assign out_psum_45 = reg_psum_63_45;
assign out_psum_46 = reg_psum_63_46;
assign out_psum_47 = reg_psum_63_47;
assign out_psum_48 = reg_psum_63_48;
assign out_psum_49 = reg_psum_63_49;
assign out_psum_50 = reg_psum_63_50;
assign out_psum_51 = reg_psum_63_51;
assign out_psum_52 = reg_psum_63_52;
assign out_psum_53 = reg_psum_63_53;
assign out_psum_54 = reg_psum_63_54;
assign out_psum_55 = reg_psum_63_55;
assign out_psum_56 = reg_psum_63_56;
assign out_psum_57 = reg_psum_63_57;
assign out_psum_58 = reg_psum_63_58;
assign out_psum_59 = reg_psum_63_59;
assign out_psum_60 = reg_psum_63_60;
assign out_psum_61 = reg_psum_63_61;
assign out_psum_62 = reg_psum_63_62;
assign out_psum_63 = reg_psum_63_63;
endmodule