`include "/home/wzc/master_project/verilog/systolic_array/PE.v"
module SA32(rst, clk, weight_en, in_weight_0, in_psum_0, in_weight_1, in_psum_1, in_weight_2, in_psum_2, in_weight_3, in_psum_3, in_weight_4, in_psum_4, in_weight_5, in_psum_5, in_weight_6, in_psum_6, in_weight_7, in_psum_7, in_weight_8, in_psum_8, in_weight_9, in_psum_9, in_weight_10, in_psum_10, in_weight_11, in_psum_11, in_weight_12, in_psum_12, in_weight_13, in_psum_13, in_weight_14, in_psum_14, in_weight_15, in_psum_15, in_weight_16, in_psum_16, in_weight_17, in_psum_17, in_weight_18, in_psum_18, in_weight_19, in_psum_19, in_weight_20, in_psum_20, in_weight_21, in_psum_21, in_weight_22, in_psum_22, in_weight_23, in_psum_23, in_weight_24, in_psum_24, in_weight_25, in_psum_25, in_weight_26, in_psum_26, in_weight_27, in_psum_27, in_weight_28, in_psum_28, in_weight_29, in_psum_29, in_weight_30, in_psum_30, in_weight_31, in_psum_31
, in_activation_0, in_activation_1, in_activation_2, in_activation_3, in_activation_4, in_activation_5, in_activation_6, in_activation_7, in_activation_8, in_activation_9, in_activation_10, in_activation_11, in_activation_12, in_activation_13, in_activation_14, in_activation_15, in_activation_16, in_activation_17, in_activation_18, in_activation_19, in_activation_20, in_activation_21, in_activation_22, in_activation_23, in_activation_24, in_activation_25, in_activation_26, in_activation_27, in_activation_28, in_activation_29, in_activation_30, in_activation_31
, out_psum_0, out_psum_1, out_psum_2, out_psum_3, out_psum_4, out_psum_5, out_psum_6, out_psum_7, out_psum_8, out_psum_9, out_psum_10, out_psum_11, out_psum_12, out_psum_13, out_psum_14, out_psum_15, out_psum_16, out_psum_17, out_psum_18, out_psum_19, out_psum_20, out_psum_21, out_psum_22, out_psum_23, out_psum_24, out_psum_25, out_psum_26, out_psum_27, out_psum_28, out_psum_29, out_psum_30, out_psum_31
, spare_out_psum_0, spare_out_psum_1, spare_out_psum_2, spare_out_psum_3, spare_out_psum_4, spare_out_psum_5, spare_out_psum_6, spare_out_psum_7, spare_out_psum_8, spare_out_psum_9, spare_out_psum_10, spare_out_psum_11, spare_out_psum_12, spare_out_psum_13, spare_out_psum_14, spare_out_psum_15, spare_out_psum_16, spare_out_psum_17, spare_out_psum_18, spare_out_psum_19, spare_out_psum_20, spare_out_psum_21, spare_out_psum_22, spare_out_psum_23, spare_out_psum_24, spare_out_psum_25, spare_out_psum_26, spare_out_psum_27, spare_out_psum_28, spare_out_psum_29, spare_out_psum_30, spare_out_psum_31);

input weight_en;
input clk,rst;
input signed[15:0]   in_weight_0;
input signed[15:0]   in_psum_0;
input signed[15:0]   in_weight_1;
input signed[15:0]   in_psum_1;
input signed[15:0]   in_weight_2;
input signed[15:0]   in_psum_2;
input signed[15:0]   in_weight_3;
input signed[15:0]   in_psum_3;
input signed[15:0]   in_weight_4;
input signed[15:0]   in_psum_4;
input signed[15:0]   in_weight_5;
input signed[15:0]   in_psum_5;
input signed[15:0]   in_weight_6;
input signed[15:0]   in_psum_6;
input signed[15:0]   in_weight_7;
input signed[15:0]   in_psum_7;
input signed[15:0]   in_weight_8;
input signed[15:0]   in_psum_8;
input signed[15:0]   in_weight_9;
input signed[15:0]   in_psum_9;
input signed[15:0]   in_weight_10;
input signed[15:0]   in_psum_10;
input signed[15:0]   in_weight_11;
input signed[15:0]   in_psum_11;
input signed[15:0]   in_weight_12;
input signed[15:0]   in_psum_12;
input signed[15:0]   in_weight_13;
input signed[15:0]   in_psum_13;
input signed[15:0]   in_weight_14;
input signed[15:0]   in_psum_14;
input signed[15:0]   in_weight_15;
input signed[15:0]   in_psum_15;
input signed[15:0]   in_weight_16;
input signed[15:0]   in_psum_16;
input signed[15:0]   in_weight_17;
input signed[15:0]   in_psum_17;
input signed[15:0]   in_weight_18;
input signed[15:0]   in_psum_18;
input signed[15:0]   in_weight_19;
input signed[15:0]   in_psum_19;
input signed[15:0]   in_weight_20;
input signed[15:0]   in_psum_20;
input signed[15:0]   in_weight_21;
input signed[15:0]   in_psum_21;
input signed[15:0]   in_weight_22;
input signed[15:0]   in_psum_22;
input signed[15:0]   in_weight_23;
input signed[15:0]   in_psum_23;
input signed[15:0]   in_weight_24;
input signed[15:0]   in_psum_24;
input signed[15:0]   in_weight_25;
input signed[15:0]   in_psum_25;
input signed[15:0]   in_weight_26;
input signed[15:0]   in_psum_26;
input signed[15:0]   in_weight_27;
input signed[15:0]   in_psum_27;
input signed[15:0]   in_weight_28;
input signed[15:0]   in_psum_28;
input signed[15:0]   in_weight_29;
input signed[15:0]   in_psum_29;
input signed[15:0]   in_weight_30;
input signed[15:0]   in_psum_30;
input signed[15:0]   in_weight_31;
input signed[15:0]   in_psum_31;
input signed[15:0]   in_activation_0;
input signed[15:0]   in_activation_1;
input signed[15:0]   in_activation_2;
input signed[15:0]   in_activation_3;
input signed[15:0]   in_activation_4;
input signed[15:0]   in_activation_5;
input signed[15:0]   in_activation_6;
input signed[15:0]   in_activation_7;
input signed[15:0]   in_activation_8;
input signed[15:0]   in_activation_9;
input signed[15:0]   in_activation_10;
input signed[15:0]   in_activation_11;
input signed[15:0]   in_activation_12;
input signed[15:0]   in_activation_13;
input signed[15:0]   in_activation_14;
input signed[15:0]   in_activation_15;
input signed[15:0]   in_activation_16;
input signed[15:0]   in_activation_17;
input signed[15:0]   in_activation_18;
input signed[15:0]   in_activation_19;
input signed[15:0]   in_activation_20;
input signed[15:0]   in_activation_21;
input signed[15:0]   in_activation_22;
input signed[15:0]   in_activation_23;
input signed[15:0]   in_activation_24;
input signed[15:0]   in_activation_25;
input signed[15:0]   in_activation_26;
input signed[15:0]   in_activation_27;
input signed[15:0]   in_activation_28;
input signed[15:0]   in_activation_29;
input signed[15:0]   in_activation_30;
input signed[15:0]   in_activation_31;
output signed[15:0]   out_psum_0;
output signed[15:0]   out_psum_1;
output signed[15:0]   out_psum_2;
output signed[15:0]   out_psum_3;
output signed[15:0]   out_psum_4;
output signed[15:0]   out_psum_5;
output signed[15:0]   out_psum_6;
output signed[15:0]   out_psum_7;
output signed[15:0]   out_psum_8;
output signed[15:0]   out_psum_9;
output signed[15:0]   out_psum_10;
output signed[15:0]   out_psum_11;
output signed[15:0]   out_psum_12;
output signed[15:0]   out_psum_13;
output signed[15:0]   out_psum_14;
output signed[15:0]   out_psum_15;
output signed[15:0]   out_psum_16;
output signed[15:0]   out_psum_17;
output signed[15:0]   out_psum_18;
output signed[15:0]   out_psum_19;
output signed[15:0]   out_psum_20;
output signed[15:0]   out_psum_21;
output signed[15:0]   out_psum_22;
output signed[15:0]   out_psum_23;
output signed[15:0]   out_psum_24;
output signed[15:0]   out_psum_25;
output signed[15:0]   out_psum_26;
output signed[15:0]   out_psum_27;
output signed[15:0]   out_psum_28;
output signed[15:0]   out_psum_29;
output signed[15:0]   out_psum_30;
output signed[15:0]   out_psum_31;
wire signed[31:0] attempt_0;
wire signed[31:0] attempt_1;
wire signed[31:0] attempt_2;
wire signed[31:0] attempt_3;
wire signed[31:0] attempt_4;
wire signed[31:0] attempt_5;
wire signed[31:0] attempt_6;
wire signed[31:0] attempt_7;
wire signed[31:0] attempt_8;
wire signed[31:0] attempt_9;
wire signed[31:0] attempt_10;
wire signed[31:0] attempt_11;
wire signed[31:0] attempt_12;
wire signed[31:0] attempt_13;
wire signed[31:0] attempt_14;
wire signed[31:0] attempt_15;
wire signed[31:0] attempt_16;
wire signed[31:0] attempt_17;
wire signed[31:0] attempt_18;
wire signed[31:0] attempt_19;
wire signed[31:0] attempt_20;
wire signed[31:0] attempt_21;
wire signed[31:0] attempt_22;
wire signed[31:0] attempt_23;
wire signed[31:0] attempt_24;
wire signed[31:0] attempt_25;
wire signed[31:0] attempt_26;
wire signed[31:0] attempt_27;
wire signed[31:0] attempt_28;
wire signed[31:0] attempt_29;
wire signed[31:0] attempt_30;
wire signed[31:0] attempt_31;
wire signed[15:0]    reg_activation_0_0;
wire signed[15:0]    reg_activation_0_1;
wire signed[15:0]    reg_activation_0_2;
wire signed[15:0]    reg_activation_0_3;
wire signed[15:0]    reg_activation_0_4;
wire signed[15:0]    reg_activation_0_5;
wire signed[15:0]    reg_activation_0_6;
wire signed[15:0]    reg_activation_0_7;
wire signed[15:0]    reg_activation_0_8;
wire signed[15:0]    reg_activation_0_9;
wire signed[15:0]    reg_activation_0_10;
wire signed[15:0]    reg_activation_0_11;
wire signed[15:0]    reg_activation_0_12;
wire signed[15:0]    reg_activation_0_13;
wire signed[15:0]    reg_activation_0_14;
wire signed[15:0]    reg_activation_0_15;
wire signed[15:0]    reg_activation_0_16;
wire signed[15:0]    reg_activation_0_17;
wire signed[15:0]    reg_activation_0_18;
wire signed[15:0]    reg_activation_0_19;
wire signed[15:0]    reg_activation_0_20;
wire signed[15:0]    reg_activation_0_21;
wire signed[15:0]    reg_activation_0_22;
wire signed[15:0]    reg_activation_0_23;
wire signed[15:0]    reg_activation_0_24;
wire signed[15:0]    reg_activation_0_25;
wire signed[15:0]    reg_activation_0_26;
wire signed[15:0]    reg_activation_0_27;
wire signed[15:0]    reg_activation_0_28;
wire signed[15:0]    reg_activation_0_29;
wire signed[15:0]    reg_activation_0_30;
wire signed[15:0]    reg_activation_0_31;
wire signed[15:0]    reg_activation_1_0;
wire signed[15:0]    reg_activation_1_1;
wire signed[15:0]    reg_activation_1_2;
wire signed[15:0]    reg_activation_1_3;
wire signed[15:0]    reg_activation_1_4;
wire signed[15:0]    reg_activation_1_5;
wire signed[15:0]    reg_activation_1_6;
wire signed[15:0]    reg_activation_1_7;
wire signed[15:0]    reg_activation_1_8;
wire signed[15:0]    reg_activation_1_9;
wire signed[15:0]    reg_activation_1_10;
wire signed[15:0]    reg_activation_1_11;
wire signed[15:0]    reg_activation_1_12;
wire signed[15:0]    reg_activation_1_13;
wire signed[15:0]    reg_activation_1_14;
wire signed[15:0]    reg_activation_1_15;
wire signed[15:0]    reg_activation_1_16;
wire signed[15:0]    reg_activation_1_17;
wire signed[15:0]    reg_activation_1_18;
wire signed[15:0]    reg_activation_1_19;
wire signed[15:0]    reg_activation_1_20;
wire signed[15:0]    reg_activation_1_21;
wire signed[15:0]    reg_activation_1_22;
wire signed[15:0]    reg_activation_1_23;
wire signed[15:0]    reg_activation_1_24;
wire signed[15:0]    reg_activation_1_25;
wire signed[15:0]    reg_activation_1_26;
wire signed[15:0]    reg_activation_1_27;
wire signed[15:0]    reg_activation_1_28;
wire signed[15:0]    reg_activation_1_29;
wire signed[15:0]    reg_activation_1_30;
wire signed[15:0]    reg_activation_1_31;
wire signed[15:0]    reg_activation_2_0;
wire signed[15:0]    reg_activation_2_1;
wire signed[15:0]    reg_activation_2_2;
wire signed[15:0]    reg_activation_2_3;
wire signed[15:0]    reg_activation_2_4;
wire signed[15:0]    reg_activation_2_5;
wire signed[15:0]    reg_activation_2_6;
wire signed[15:0]    reg_activation_2_7;
wire signed[15:0]    reg_activation_2_8;
wire signed[15:0]    reg_activation_2_9;
wire signed[15:0]    reg_activation_2_10;
wire signed[15:0]    reg_activation_2_11;
wire signed[15:0]    reg_activation_2_12;
wire signed[15:0]    reg_activation_2_13;
wire signed[15:0]    reg_activation_2_14;
wire signed[15:0]    reg_activation_2_15;
wire signed[15:0]    reg_activation_2_16;
wire signed[15:0]    reg_activation_2_17;
wire signed[15:0]    reg_activation_2_18;
wire signed[15:0]    reg_activation_2_19;
wire signed[15:0]    reg_activation_2_20;
wire signed[15:0]    reg_activation_2_21;
wire signed[15:0]    reg_activation_2_22;
wire signed[15:0]    reg_activation_2_23;
wire signed[15:0]    reg_activation_2_24;
wire signed[15:0]    reg_activation_2_25;
wire signed[15:0]    reg_activation_2_26;
wire signed[15:0]    reg_activation_2_27;
wire signed[15:0]    reg_activation_2_28;
wire signed[15:0]    reg_activation_2_29;
wire signed[15:0]    reg_activation_2_30;
wire signed[15:0]    reg_activation_2_31;
wire signed[15:0]    reg_activation_3_0;
wire signed[15:0]    reg_activation_3_1;
wire signed[15:0]    reg_activation_3_2;
wire signed[15:0]    reg_activation_3_3;
wire signed[15:0]    reg_activation_3_4;
wire signed[15:0]    reg_activation_3_5;
wire signed[15:0]    reg_activation_3_6;
wire signed[15:0]    reg_activation_3_7;
wire signed[15:0]    reg_activation_3_8;
wire signed[15:0]    reg_activation_3_9;
wire signed[15:0]    reg_activation_3_10;
wire signed[15:0]    reg_activation_3_11;
wire signed[15:0]    reg_activation_3_12;
wire signed[15:0]    reg_activation_3_13;
wire signed[15:0]    reg_activation_3_14;
wire signed[15:0]    reg_activation_3_15;
wire signed[15:0]    reg_activation_3_16;
wire signed[15:0]    reg_activation_3_17;
wire signed[15:0]    reg_activation_3_18;
wire signed[15:0]    reg_activation_3_19;
wire signed[15:0]    reg_activation_3_20;
wire signed[15:0]    reg_activation_3_21;
wire signed[15:0]    reg_activation_3_22;
wire signed[15:0]    reg_activation_3_23;
wire signed[15:0]    reg_activation_3_24;
wire signed[15:0]    reg_activation_3_25;
wire signed[15:0]    reg_activation_3_26;
wire signed[15:0]    reg_activation_3_27;
wire signed[15:0]    reg_activation_3_28;
wire signed[15:0]    reg_activation_3_29;
wire signed[15:0]    reg_activation_3_30;
wire signed[15:0]    reg_activation_3_31;
wire signed[15:0]    reg_activation_4_0;
wire signed[15:0]    reg_activation_4_1;
wire signed[15:0]    reg_activation_4_2;
wire signed[15:0]    reg_activation_4_3;
wire signed[15:0]    reg_activation_4_4;
wire signed[15:0]    reg_activation_4_5;
wire signed[15:0]    reg_activation_4_6;
wire signed[15:0]    reg_activation_4_7;
wire signed[15:0]    reg_activation_4_8;
wire signed[15:0]    reg_activation_4_9;
wire signed[15:0]    reg_activation_4_10;
wire signed[15:0]    reg_activation_4_11;
wire signed[15:0]    reg_activation_4_12;
wire signed[15:0]    reg_activation_4_13;
wire signed[15:0]    reg_activation_4_14;
wire signed[15:0]    reg_activation_4_15;
wire signed[15:0]    reg_activation_4_16;
wire signed[15:0]    reg_activation_4_17;
wire signed[15:0]    reg_activation_4_18;
wire signed[15:0]    reg_activation_4_19;
wire signed[15:0]    reg_activation_4_20;
wire signed[15:0]    reg_activation_4_21;
wire signed[15:0]    reg_activation_4_22;
wire signed[15:0]    reg_activation_4_23;
wire signed[15:0]    reg_activation_4_24;
wire signed[15:0]    reg_activation_4_25;
wire signed[15:0]    reg_activation_4_26;
wire signed[15:0]    reg_activation_4_27;
wire signed[15:0]    reg_activation_4_28;
wire signed[15:0]    reg_activation_4_29;
wire signed[15:0]    reg_activation_4_30;
wire signed[15:0]    reg_activation_4_31;
wire signed[15:0]    reg_activation_5_0;
wire signed[15:0]    reg_activation_5_1;
wire signed[15:0]    reg_activation_5_2;
wire signed[15:0]    reg_activation_5_3;
wire signed[15:0]    reg_activation_5_4;
wire signed[15:0]    reg_activation_5_5;
wire signed[15:0]    reg_activation_5_6;
wire signed[15:0]    reg_activation_5_7;
wire signed[15:0]    reg_activation_5_8;
wire signed[15:0]    reg_activation_5_9;
wire signed[15:0]    reg_activation_5_10;
wire signed[15:0]    reg_activation_5_11;
wire signed[15:0]    reg_activation_5_12;
wire signed[15:0]    reg_activation_5_13;
wire signed[15:0]    reg_activation_5_14;
wire signed[15:0]    reg_activation_5_15;
wire signed[15:0]    reg_activation_5_16;
wire signed[15:0]    reg_activation_5_17;
wire signed[15:0]    reg_activation_5_18;
wire signed[15:0]    reg_activation_5_19;
wire signed[15:0]    reg_activation_5_20;
wire signed[15:0]    reg_activation_5_21;
wire signed[15:0]    reg_activation_5_22;
wire signed[15:0]    reg_activation_5_23;
wire signed[15:0]    reg_activation_5_24;
wire signed[15:0]    reg_activation_5_25;
wire signed[15:0]    reg_activation_5_26;
wire signed[15:0]    reg_activation_5_27;
wire signed[15:0]    reg_activation_5_28;
wire signed[15:0]    reg_activation_5_29;
wire signed[15:0]    reg_activation_5_30;
wire signed[15:0]    reg_activation_5_31;
wire signed[15:0]    reg_activation_6_0;
wire signed[15:0]    reg_activation_6_1;
wire signed[15:0]    reg_activation_6_2;
wire signed[15:0]    reg_activation_6_3;
wire signed[15:0]    reg_activation_6_4;
wire signed[15:0]    reg_activation_6_5;
wire signed[15:0]    reg_activation_6_6;
wire signed[15:0]    reg_activation_6_7;
wire signed[15:0]    reg_activation_6_8;
wire signed[15:0]    reg_activation_6_9;
wire signed[15:0]    reg_activation_6_10;
wire signed[15:0]    reg_activation_6_11;
wire signed[15:0]    reg_activation_6_12;
wire signed[15:0]    reg_activation_6_13;
wire signed[15:0]    reg_activation_6_14;
wire signed[15:0]    reg_activation_6_15;
wire signed[15:0]    reg_activation_6_16;
wire signed[15:0]    reg_activation_6_17;
wire signed[15:0]    reg_activation_6_18;
wire signed[15:0]    reg_activation_6_19;
wire signed[15:0]    reg_activation_6_20;
wire signed[15:0]    reg_activation_6_21;
wire signed[15:0]    reg_activation_6_22;
wire signed[15:0]    reg_activation_6_23;
wire signed[15:0]    reg_activation_6_24;
wire signed[15:0]    reg_activation_6_25;
wire signed[15:0]    reg_activation_6_26;
wire signed[15:0]    reg_activation_6_27;
wire signed[15:0]    reg_activation_6_28;
wire signed[15:0]    reg_activation_6_29;
wire signed[15:0]    reg_activation_6_30;
wire signed[15:0]    reg_activation_6_31;
wire signed[15:0]    reg_activation_7_0;
wire signed[15:0]    reg_activation_7_1;
wire signed[15:0]    reg_activation_7_2;
wire signed[15:0]    reg_activation_7_3;
wire signed[15:0]    reg_activation_7_4;
wire signed[15:0]    reg_activation_7_5;
wire signed[15:0]    reg_activation_7_6;
wire signed[15:0]    reg_activation_7_7;
wire signed[15:0]    reg_activation_7_8;
wire signed[15:0]    reg_activation_7_9;
wire signed[15:0]    reg_activation_7_10;
wire signed[15:0]    reg_activation_7_11;
wire signed[15:0]    reg_activation_7_12;
wire signed[15:0]    reg_activation_7_13;
wire signed[15:0]    reg_activation_7_14;
wire signed[15:0]    reg_activation_7_15;
wire signed[15:0]    reg_activation_7_16;
wire signed[15:0]    reg_activation_7_17;
wire signed[15:0]    reg_activation_7_18;
wire signed[15:0]    reg_activation_7_19;
wire signed[15:0]    reg_activation_7_20;
wire signed[15:0]    reg_activation_7_21;
wire signed[15:0]    reg_activation_7_22;
wire signed[15:0]    reg_activation_7_23;
wire signed[15:0]    reg_activation_7_24;
wire signed[15:0]    reg_activation_7_25;
wire signed[15:0]    reg_activation_7_26;
wire signed[15:0]    reg_activation_7_27;
wire signed[15:0]    reg_activation_7_28;
wire signed[15:0]    reg_activation_7_29;
wire signed[15:0]    reg_activation_7_30;
wire signed[15:0]    reg_activation_7_31;
wire signed[15:0]    reg_activation_8_0;
wire signed[15:0]    reg_activation_8_1;
wire signed[15:0]    reg_activation_8_2;
wire signed[15:0]    reg_activation_8_3;
wire signed[15:0]    reg_activation_8_4;
wire signed[15:0]    reg_activation_8_5;
wire signed[15:0]    reg_activation_8_6;
wire signed[15:0]    reg_activation_8_7;
wire signed[15:0]    reg_activation_8_8;
wire signed[15:0]    reg_activation_8_9;
wire signed[15:0]    reg_activation_8_10;
wire signed[15:0]    reg_activation_8_11;
wire signed[15:0]    reg_activation_8_12;
wire signed[15:0]    reg_activation_8_13;
wire signed[15:0]    reg_activation_8_14;
wire signed[15:0]    reg_activation_8_15;
wire signed[15:0]    reg_activation_8_16;
wire signed[15:0]    reg_activation_8_17;
wire signed[15:0]    reg_activation_8_18;
wire signed[15:0]    reg_activation_8_19;
wire signed[15:0]    reg_activation_8_20;
wire signed[15:0]    reg_activation_8_21;
wire signed[15:0]    reg_activation_8_22;
wire signed[15:0]    reg_activation_8_23;
wire signed[15:0]    reg_activation_8_24;
wire signed[15:0]    reg_activation_8_25;
wire signed[15:0]    reg_activation_8_26;
wire signed[15:0]    reg_activation_8_27;
wire signed[15:0]    reg_activation_8_28;
wire signed[15:0]    reg_activation_8_29;
wire signed[15:0]    reg_activation_8_30;
wire signed[15:0]    reg_activation_8_31;
wire signed[15:0]    reg_activation_9_0;
wire signed[15:0]    reg_activation_9_1;
wire signed[15:0]    reg_activation_9_2;
wire signed[15:0]    reg_activation_9_3;
wire signed[15:0]    reg_activation_9_4;
wire signed[15:0]    reg_activation_9_5;
wire signed[15:0]    reg_activation_9_6;
wire signed[15:0]    reg_activation_9_7;
wire signed[15:0]    reg_activation_9_8;
wire signed[15:0]    reg_activation_9_9;
wire signed[15:0]    reg_activation_9_10;
wire signed[15:0]    reg_activation_9_11;
wire signed[15:0]    reg_activation_9_12;
wire signed[15:0]    reg_activation_9_13;
wire signed[15:0]    reg_activation_9_14;
wire signed[15:0]    reg_activation_9_15;
wire signed[15:0]    reg_activation_9_16;
wire signed[15:0]    reg_activation_9_17;
wire signed[15:0]    reg_activation_9_18;
wire signed[15:0]    reg_activation_9_19;
wire signed[15:0]    reg_activation_9_20;
wire signed[15:0]    reg_activation_9_21;
wire signed[15:0]    reg_activation_9_22;
wire signed[15:0]    reg_activation_9_23;
wire signed[15:0]    reg_activation_9_24;
wire signed[15:0]    reg_activation_9_25;
wire signed[15:0]    reg_activation_9_26;
wire signed[15:0]    reg_activation_9_27;
wire signed[15:0]    reg_activation_9_28;
wire signed[15:0]    reg_activation_9_29;
wire signed[15:0]    reg_activation_9_30;
wire signed[15:0]    reg_activation_9_31;
wire signed[15:0]    reg_activation_10_0;
wire signed[15:0]    reg_activation_10_1;
wire signed[15:0]    reg_activation_10_2;
wire signed[15:0]    reg_activation_10_3;
wire signed[15:0]    reg_activation_10_4;
wire signed[15:0]    reg_activation_10_5;
wire signed[15:0]    reg_activation_10_6;
wire signed[15:0]    reg_activation_10_7;
wire signed[15:0]    reg_activation_10_8;
wire signed[15:0]    reg_activation_10_9;
wire signed[15:0]    reg_activation_10_10;
wire signed[15:0]    reg_activation_10_11;
wire signed[15:0]    reg_activation_10_12;
wire signed[15:0]    reg_activation_10_13;
wire signed[15:0]    reg_activation_10_14;
wire signed[15:0]    reg_activation_10_15;
wire signed[15:0]    reg_activation_10_16;
wire signed[15:0]    reg_activation_10_17;
wire signed[15:0]    reg_activation_10_18;
wire signed[15:0]    reg_activation_10_19;
wire signed[15:0]    reg_activation_10_20;
wire signed[15:0]    reg_activation_10_21;
wire signed[15:0]    reg_activation_10_22;
wire signed[15:0]    reg_activation_10_23;
wire signed[15:0]    reg_activation_10_24;
wire signed[15:0]    reg_activation_10_25;
wire signed[15:0]    reg_activation_10_26;
wire signed[15:0]    reg_activation_10_27;
wire signed[15:0]    reg_activation_10_28;
wire signed[15:0]    reg_activation_10_29;
wire signed[15:0]    reg_activation_10_30;
wire signed[15:0]    reg_activation_10_31;
wire signed[15:0]    reg_activation_11_0;
wire signed[15:0]    reg_activation_11_1;
wire signed[15:0]    reg_activation_11_2;
wire signed[15:0]    reg_activation_11_3;
wire signed[15:0]    reg_activation_11_4;
wire signed[15:0]    reg_activation_11_5;
wire signed[15:0]    reg_activation_11_6;
wire signed[15:0]    reg_activation_11_7;
wire signed[15:0]    reg_activation_11_8;
wire signed[15:0]    reg_activation_11_9;
wire signed[15:0]    reg_activation_11_10;
wire signed[15:0]    reg_activation_11_11;
wire signed[15:0]    reg_activation_11_12;
wire signed[15:0]    reg_activation_11_13;
wire signed[15:0]    reg_activation_11_14;
wire signed[15:0]    reg_activation_11_15;
wire signed[15:0]    reg_activation_11_16;
wire signed[15:0]    reg_activation_11_17;
wire signed[15:0]    reg_activation_11_18;
wire signed[15:0]    reg_activation_11_19;
wire signed[15:0]    reg_activation_11_20;
wire signed[15:0]    reg_activation_11_21;
wire signed[15:0]    reg_activation_11_22;
wire signed[15:0]    reg_activation_11_23;
wire signed[15:0]    reg_activation_11_24;
wire signed[15:0]    reg_activation_11_25;
wire signed[15:0]    reg_activation_11_26;
wire signed[15:0]    reg_activation_11_27;
wire signed[15:0]    reg_activation_11_28;
wire signed[15:0]    reg_activation_11_29;
wire signed[15:0]    reg_activation_11_30;
wire signed[15:0]    reg_activation_11_31;
wire signed[15:0]    reg_activation_12_0;
wire signed[15:0]    reg_activation_12_1;
wire signed[15:0]    reg_activation_12_2;
wire signed[15:0]    reg_activation_12_3;
wire signed[15:0]    reg_activation_12_4;
wire signed[15:0]    reg_activation_12_5;
wire signed[15:0]    reg_activation_12_6;
wire signed[15:0]    reg_activation_12_7;
wire signed[15:0]    reg_activation_12_8;
wire signed[15:0]    reg_activation_12_9;
wire signed[15:0]    reg_activation_12_10;
wire signed[15:0]    reg_activation_12_11;
wire signed[15:0]    reg_activation_12_12;
wire signed[15:0]    reg_activation_12_13;
wire signed[15:0]    reg_activation_12_14;
wire signed[15:0]    reg_activation_12_15;
wire signed[15:0]    reg_activation_12_16;
wire signed[15:0]    reg_activation_12_17;
wire signed[15:0]    reg_activation_12_18;
wire signed[15:0]    reg_activation_12_19;
wire signed[15:0]    reg_activation_12_20;
wire signed[15:0]    reg_activation_12_21;
wire signed[15:0]    reg_activation_12_22;
wire signed[15:0]    reg_activation_12_23;
wire signed[15:0]    reg_activation_12_24;
wire signed[15:0]    reg_activation_12_25;
wire signed[15:0]    reg_activation_12_26;
wire signed[15:0]    reg_activation_12_27;
wire signed[15:0]    reg_activation_12_28;
wire signed[15:0]    reg_activation_12_29;
wire signed[15:0]    reg_activation_12_30;
wire signed[15:0]    reg_activation_12_31;
wire signed[15:0]    reg_activation_13_0;
wire signed[15:0]    reg_activation_13_1;
wire signed[15:0]    reg_activation_13_2;
wire signed[15:0]    reg_activation_13_3;
wire signed[15:0]    reg_activation_13_4;
wire signed[15:0]    reg_activation_13_5;
wire signed[15:0]    reg_activation_13_6;
wire signed[15:0]    reg_activation_13_7;
wire signed[15:0]    reg_activation_13_8;
wire signed[15:0]    reg_activation_13_9;
wire signed[15:0]    reg_activation_13_10;
wire signed[15:0]    reg_activation_13_11;
wire signed[15:0]    reg_activation_13_12;
wire signed[15:0]    reg_activation_13_13;
wire signed[15:0]    reg_activation_13_14;
wire signed[15:0]    reg_activation_13_15;
wire signed[15:0]    reg_activation_13_16;
wire signed[15:0]    reg_activation_13_17;
wire signed[15:0]    reg_activation_13_18;
wire signed[15:0]    reg_activation_13_19;
wire signed[15:0]    reg_activation_13_20;
wire signed[15:0]    reg_activation_13_21;
wire signed[15:0]    reg_activation_13_22;
wire signed[15:0]    reg_activation_13_23;
wire signed[15:0]    reg_activation_13_24;
wire signed[15:0]    reg_activation_13_25;
wire signed[15:0]    reg_activation_13_26;
wire signed[15:0]    reg_activation_13_27;
wire signed[15:0]    reg_activation_13_28;
wire signed[15:0]    reg_activation_13_29;
wire signed[15:0]    reg_activation_13_30;
wire signed[15:0]    reg_activation_13_31;
wire signed[15:0]    reg_activation_14_0;
wire signed[15:0]    reg_activation_14_1;
wire signed[15:0]    reg_activation_14_2;
wire signed[15:0]    reg_activation_14_3;
wire signed[15:0]    reg_activation_14_4;
wire signed[15:0]    reg_activation_14_5;
wire signed[15:0]    reg_activation_14_6;
wire signed[15:0]    reg_activation_14_7;
wire signed[15:0]    reg_activation_14_8;
wire signed[15:0]    reg_activation_14_9;
wire signed[15:0]    reg_activation_14_10;
wire signed[15:0]    reg_activation_14_11;
wire signed[15:0]    reg_activation_14_12;
wire signed[15:0]    reg_activation_14_13;
wire signed[15:0]    reg_activation_14_14;
wire signed[15:0]    reg_activation_14_15;
wire signed[15:0]    reg_activation_14_16;
wire signed[15:0]    reg_activation_14_17;
wire signed[15:0]    reg_activation_14_18;
wire signed[15:0]    reg_activation_14_19;
wire signed[15:0]    reg_activation_14_20;
wire signed[15:0]    reg_activation_14_21;
wire signed[15:0]    reg_activation_14_22;
wire signed[15:0]    reg_activation_14_23;
wire signed[15:0]    reg_activation_14_24;
wire signed[15:0]    reg_activation_14_25;
wire signed[15:0]    reg_activation_14_26;
wire signed[15:0]    reg_activation_14_27;
wire signed[15:0]    reg_activation_14_28;
wire signed[15:0]    reg_activation_14_29;
wire signed[15:0]    reg_activation_14_30;
wire signed[15:0]    reg_activation_14_31;
wire signed[15:0]    reg_activation_15_0;
wire signed[15:0]    reg_activation_15_1;
wire signed[15:0]    reg_activation_15_2;
wire signed[15:0]    reg_activation_15_3;
wire signed[15:0]    reg_activation_15_4;
wire signed[15:0]    reg_activation_15_5;
wire signed[15:0]    reg_activation_15_6;
wire signed[15:0]    reg_activation_15_7;
wire signed[15:0]    reg_activation_15_8;
wire signed[15:0]    reg_activation_15_9;
wire signed[15:0]    reg_activation_15_10;
wire signed[15:0]    reg_activation_15_11;
wire signed[15:0]    reg_activation_15_12;
wire signed[15:0]    reg_activation_15_13;
wire signed[15:0]    reg_activation_15_14;
wire signed[15:0]    reg_activation_15_15;
wire signed[15:0]    reg_activation_15_16;
wire signed[15:0]    reg_activation_15_17;
wire signed[15:0]    reg_activation_15_18;
wire signed[15:0]    reg_activation_15_19;
wire signed[15:0]    reg_activation_15_20;
wire signed[15:0]    reg_activation_15_21;
wire signed[15:0]    reg_activation_15_22;
wire signed[15:0]    reg_activation_15_23;
wire signed[15:0]    reg_activation_15_24;
wire signed[15:0]    reg_activation_15_25;
wire signed[15:0]    reg_activation_15_26;
wire signed[15:0]    reg_activation_15_27;
wire signed[15:0]    reg_activation_15_28;
wire signed[15:0]    reg_activation_15_29;
wire signed[15:0]    reg_activation_15_30;
wire signed[15:0]    reg_activation_15_31;
wire signed[15:0]    reg_activation_16_0;
wire signed[15:0]    reg_activation_16_1;
wire signed[15:0]    reg_activation_16_2;
wire signed[15:0]    reg_activation_16_3;
wire signed[15:0]    reg_activation_16_4;
wire signed[15:0]    reg_activation_16_5;
wire signed[15:0]    reg_activation_16_6;
wire signed[15:0]    reg_activation_16_7;
wire signed[15:0]    reg_activation_16_8;
wire signed[15:0]    reg_activation_16_9;
wire signed[15:0]    reg_activation_16_10;
wire signed[15:0]    reg_activation_16_11;
wire signed[15:0]    reg_activation_16_12;
wire signed[15:0]    reg_activation_16_13;
wire signed[15:0]    reg_activation_16_14;
wire signed[15:0]    reg_activation_16_15;
wire signed[15:0]    reg_activation_16_16;
wire signed[15:0]    reg_activation_16_17;
wire signed[15:0]    reg_activation_16_18;
wire signed[15:0]    reg_activation_16_19;
wire signed[15:0]    reg_activation_16_20;
wire signed[15:0]    reg_activation_16_21;
wire signed[15:0]    reg_activation_16_22;
wire signed[15:0]    reg_activation_16_23;
wire signed[15:0]    reg_activation_16_24;
wire signed[15:0]    reg_activation_16_25;
wire signed[15:0]    reg_activation_16_26;
wire signed[15:0]    reg_activation_16_27;
wire signed[15:0]    reg_activation_16_28;
wire signed[15:0]    reg_activation_16_29;
wire signed[15:0]    reg_activation_16_30;
wire signed[15:0]    reg_activation_16_31;
wire signed[15:0]    reg_activation_17_0;
wire signed[15:0]    reg_activation_17_1;
wire signed[15:0]    reg_activation_17_2;
wire signed[15:0]    reg_activation_17_3;
wire signed[15:0]    reg_activation_17_4;
wire signed[15:0]    reg_activation_17_5;
wire signed[15:0]    reg_activation_17_6;
wire signed[15:0]    reg_activation_17_7;
wire signed[15:0]    reg_activation_17_8;
wire signed[15:0]    reg_activation_17_9;
wire signed[15:0]    reg_activation_17_10;
wire signed[15:0]    reg_activation_17_11;
wire signed[15:0]    reg_activation_17_12;
wire signed[15:0]    reg_activation_17_13;
wire signed[15:0]    reg_activation_17_14;
wire signed[15:0]    reg_activation_17_15;
wire signed[15:0]    reg_activation_17_16;
wire signed[15:0]    reg_activation_17_17;
wire signed[15:0]    reg_activation_17_18;
wire signed[15:0]    reg_activation_17_19;
wire signed[15:0]    reg_activation_17_20;
wire signed[15:0]    reg_activation_17_21;
wire signed[15:0]    reg_activation_17_22;
wire signed[15:0]    reg_activation_17_23;
wire signed[15:0]    reg_activation_17_24;
wire signed[15:0]    reg_activation_17_25;
wire signed[15:0]    reg_activation_17_26;
wire signed[15:0]    reg_activation_17_27;
wire signed[15:0]    reg_activation_17_28;
wire signed[15:0]    reg_activation_17_29;
wire signed[15:0]    reg_activation_17_30;
wire signed[15:0]    reg_activation_17_31;
wire signed[15:0]    reg_activation_18_0;
wire signed[15:0]    reg_activation_18_1;
wire signed[15:0]    reg_activation_18_2;
wire signed[15:0]    reg_activation_18_3;
wire signed[15:0]    reg_activation_18_4;
wire signed[15:0]    reg_activation_18_5;
wire signed[15:0]    reg_activation_18_6;
wire signed[15:0]    reg_activation_18_7;
wire signed[15:0]    reg_activation_18_8;
wire signed[15:0]    reg_activation_18_9;
wire signed[15:0]    reg_activation_18_10;
wire signed[15:0]    reg_activation_18_11;
wire signed[15:0]    reg_activation_18_12;
wire signed[15:0]    reg_activation_18_13;
wire signed[15:0]    reg_activation_18_14;
wire signed[15:0]    reg_activation_18_15;
wire signed[15:0]    reg_activation_18_16;
wire signed[15:0]    reg_activation_18_17;
wire signed[15:0]    reg_activation_18_18;
wire signed[15:0]    reg_activation_18_19;
wire signed[15:0]    reg_activation_18_20;
wire signed[15:0]    reg_activation_18_21;
wire signed[15:0]    reg_activation_18_22;
wire signed[15:0]    reg_activation_18_23;
wire signed[15:0]    reg_activation_18_24;
wire signed[15:0]    reg_activation_18_25;
wire signed[15:0]    reg_activation_18_26;
wire signed[15:0]    reg_activation_18_27;
wire signed[15:0]    reg_activation_18_28;
wire signed[15:0]    reg_activation_18_29;
wire signed[15:0]    reg_activation_18_30;
wire signed[15:0]    reg_activation_18_31;
wire signed[15:0]    reg_activation_19_0;
wire signed[15:0]    reg_activation_19_1;
wire signed[15:0]    reg_activation_19_2;
wire signed[15:0]    reg_activation_19_3;
wire signed[15:0]    reg_activation_19_4;
wire signed[15:0]    reg_activation_19_5;
wire signed[15:0]    reg_activation_19_6;
wire signed[15:0]    reg_activation_19_7;
wire signed[15:0]    reg_activation_19_8;
wire signed[15:0]    reg_activation_19_9;
wire signed[15:0]    reg_activation_19_10;
wire signed[15:0]    reg_activation_19_11;
wire signed[15:0]    reg_activation_19_12;
wire signed[15:0]    reg_activation_19_13;
wire signed[15:0]    reg_activation_19_14;
wire signed[15:0]    reg_activation_19_15;
wire signed[15:0]    reg_activation_19_16;
wire signed[15:0]    reg_activation_19_17;
wire signed[15:0]    reg_activation_19_18;
wire signed[15:0]    reg_activation_19_19;
wire signed[15:0]    reg_activation_19_20;
wire signed[15:0]    reg_activation_19_21;
wire signed[15:0]    reg_activation_19_22;
wire signed[15:0]    reg_activation_19_23;
wire signed[15:0]    reg_activation_19_24;
wire signed[15:0]    reg_activation_19_25;
wire signed[15:0]    reg_activation_19_26;
wire signed[15:0]    reg_activation_19_27;
wire signed[15:0]    reg_activation_19_28;
wire signed[15:0]    reg_activation_19_29;
wire signed[15:0]    reg_activation_19_30;
wire signed[15:0]    reg_activation_19_31;
wire signed[15:0]    reg_activation_20_0;
wire signed[15:0]    reg_activation_20_1;
wire signed[15:0]    reg_activation_20_2;
wire signed[15:0]    reg_activation_20_3;
wire signed[15:0]    reg_activation_20_4;
wire signed[15:0]    reg_activation_20_5;
wire signed[15:0]    reg_activation_20_6;
wire signed[15:0]    reg_activation_20_7;
wire signed[15:0]    reg_activation_20_8;
wire signed[15:0]    reg_activation_20_9;
wire signed[15:0]    reg_activation_20_10;
wire signed[15:0]    reg_activation_20_11;
wire signed[15:0]    reg_activation_20_12;
wire signed[15:0]    reg_activation_20_13;
wire signed[15:0]    reg_activation_20_14;
wire signed[15:0]    reg_activation_20_15;
wire signed[15:0]    reg_activation_20_16;
wire signed[15:0]    reg_activation_20_17;
wire signed[15:0]    reg_activation_20_18;
wire signed[15:0]    reg_activation_20_19;
wire signed[15:0]    reg_activation_20_20;
wire signed[15:0]    reg_activation_20_21;
wire signed[15:0]    reg_activation_20_22;
wire signed[15:0]    reg_activation_20_23;
wire signed[15:0]    reg_activation_20_24;
wire signed[15:0]    reg_activation_20_25;
wire signed[15:0]    reg_activation_20_26;
wire signed[15:0]    reg_activation_20_27;
wire signed[15:0]    reg_activation_20_28;
wire signed[15:0]    reg_activation_20_29;
wire signed[15:0]    reg_activation_20_30;
wire signed[15:0]    reg_activation_20_31;
wire signed[15:0]    reg_activation_21_0;
wire signed[15:0]    reg_activation_21_1;
wire signed[15:0]    reg_activation_21_2;
wire signed[15:0]    reg_activation_21_3;
wire signed[15:0]    reg_activation_21_4;
wire signed[15:0]    reg_activation_21_5;
wire signed[15:0]    reg_activation_21_6;
wire signed[15:0]    reg_activation_21_7;
wire signed[15:0]    reg_activation_21_8;
wire signed[15:0]    reg_activation_21_9;
wire signed[15:0]    reg_activation_21_10;
wire signed[15:0]    reg_activation_21_11;
wire signed[15:0]    reg_activation_21_12;
wire signed[15:0]    reg_activation_21_13;
wire signed[15:0]    reg_activation_21_14;
wire signed[15:0]    reg_activation_21_15;
wire signed[15:0]    reg_activation_21_16;
wire signed[15:0]    reg_activation_21_17;
wire signed[15:0]    reg_activation_21_18;
wire signed[15:0]    reg_activation_21_19;
wire signed[15:0]    reg_activation_21_20;
wire signed[15:0]    reg_activation_21_21;
wire signed[15:0]    reg_activation_21_22;
wire signed[15:0]    reg_activation_21_23;
wire signed[15:0]    reg_activation_21_24;
wire signed[15:0]    reg_activation_21_25;
wire signed[15:0]    reg_activation_21_26;
wire signed[15:0]    reg_activation_21_27;
wire signed[15:0]    reg_activation_21_28;
wire signed[15:0]    reg_activation_21_29;
wire signed[15:0]    reg_activation_21_30;
wire signed[15:0]    reg_activation_21_31;
wire signed[15:0]    reg_activation_22_0;
wire signed[15:0]    reg_activation_22_1;
wire signed[15:0]    reg_activation_22_2;
wire signed[15:0]    reg_activation_22_3;
wire signed[15:0]    reg_activation_22_4;
wire signed[15:0]    reg_activation_22_5;
wire signed[15:0]    reg_activation_22_6;
wire signed[15:0]    reg_activation_22_7;
wire signed[15:0]    reg_activation_22_8;
wire signed[15:0]    reg_activation_22_9;
wire signed[15:0]    reg_activation_22_10;
wire signed[15:0]    reg_activation_22_11;
wire signed[15:0]    reg_activation_22_12;
wire signed[15:0]    reg_activation_22_13;
wire signed[15:0]    reg_activation_22_14;
wire signed[15:0]    reg_activation_22_15;
wire signed[15:0]    reg_activation_22_16;
wire signed[15:0]    reg_activation_22_17;
wire signed[15:0]    reg_activation_22_18;
wire signed[15:0]    reg_activation_22_19;
wire signed[15:0]    reg_activation_22_20;
wire signed[15:0]    reg_activation_22_21;
wire signed[15:0]    reg_activation_22_22;
wire signed[15:0]    reg_activation_22_23;
wire signed[15:0]    reg_activation_22_24;
wire signed[15:0]    reg_activation_22_25;
wire signed[15:0]    reg_activation_22_26;
wire signed[15:0]    reg_activation_22_27;
wire signed[15:0]    reg_activation_22_28;
wire signed[15:0]    reg_activation_22_29;
wire signed[15:0]    reg_activation_22_30;
wire signed[15:0]    reg_activation_22_31;
wire signed[15:0]    reg_activation_23_0;
wire signed[15:0]    reg_activation_23_1;
wire signed[15:0]    reg_activation_23_2;
wire signed[15:0]    reg_activation_23_3;
wire signed[15:0]    reg_activation_23_4;
wire signed[15:0]    reg_activation_23_5;
wire signed[15:0]    reg_activation_23_6;
wire signed[15:0]    reg_activation_23_7;
wire signed[15:0]    reg_activation_23_8;
wire signed[15:0]    reg_activation_23_9;
wire signed[15:0]    reg_activation_23_10;
wire signed[15:0]    reg_activation_23_11;
wire signed[15:0]    reg_activation_23_12;
wire signed[15:0]    reg_activation_23_13;
wire signed[15:0]    reg_activation_23_14;
wire signed[15:0]    reg_activation_23_15;
wire signed[15:0]    reg_activation_23_16;
wire signed[15:0]    reg_activation_23_17;
wire signed[15:0]    reg_activation_23_18;
wire signed[15:0]    reg_activation_23_19;
wire signed[15:0]    reg_activation_23_20;
wire signed[15:0]    reg_activation_23_21;
wire signed[15:0]    reg_activation_23_22;
wire signed[15:0]    reg_activation_23_23;
wire signed[15:0]    reg_activation_23_24;
wire signed[15:0]    reg_activation_23_25;
wire signed[15:0]    reg_activation_23_26;
wire signed[15:0]    reg_activation_23_27;
wire signed[15:0]    reg_activation_23_28;
wire signed[15:0]    reg_activation_23_29;
wire signed[15:0]    reg_activation_23_30;
wire signed[15:0]    reg_activation_23_31;
wire signed[15:0]    reg_activation_24_0;
wire signed[15:0]    reg_activation_24_1;
wire signed[15:0]    reg_activation_24_2;
wire signed[15:0]    reg_activation_24_3;
wire signed[15:0]    reg_activation_24_4;
wire signed[15:0]    reg_activation_24_5;
wire signed[15:0]    reg_activation_24_6;
wire signed[15:0]    reg_activation_24_7;
wire signed[15:0]    reg_activation_24_8;
wire signed[15:0]    reg_activation_24_9;
wire signed[15:0]    reg_activation_24_10;
wire signed[15:0]    reg_activation_24_11;
wire signed[15:0]    reg_activation_24_12;
wire signed[15:0]    reg_activation_24_13;
wire signed[15:0]    reg_activation_24_14;
wire signed[15:0]    reg_activation_24_15;
wire signed[15:0]    reg_activation_24_16;
wire signed[15:0]    reg_activation_24_17;
wire signed[15:0]    reg_activation_24_18;
wire signed[15:0]    reg_activation_24_19;
wire signed[15:0]    reg_activation_24_20;
wire signed[15:0]    reg_activation_24_21;
wire signed[15:0]    reg_activation_24_22;
wire signed[15:0]    reg_activation_24_23;
wire signed[15:0]    reg_activation_24_24;
wire signed[15:0]    reg_activation_24_25;
wire signed[15:0]    reg_activation_24_26;
wire signed[15:0]    reg_activation_24_27;
wire signed[15:0]    reg_activation_24_28;
wire signed[15:0]    reg_activation_24_29;
wire signed[15:0]    reg_activation_24_30;
wire signed[15:0]    reg_activation_24_31;
wire signed[15:0]    reg_activation_25_0;
wire signed[15:0]    reg_activation_25_1;
wire signed[15:0]    reg_activation_25_2;
wire signed[15:0]    reg_activation_25_3;
wire signed[15:0]    reg_activation_25_4;
wire signed[15:0]    reg_activation_25_5;
wire signed[15:0]    reg_activation_25_6;
wire signed[15:0]    reg_activation_25_7;
wire signed[15:0]    reg_activation_25_8;
wire signed[15:0]    reg_activation_25_9;
wire signed[15:0]    reg_activation_25_10;
wire signed[15:0]    reg_activation_25_11;
wire signed[15:0]    reg_activation_25_12;
wire signed[15:0]    reg_activation_25_13;
wire signed[15:0]    reg_activation_25_14;
wire signed[15:0]    reg_activation_25_15;
wire signed[15:0]    reg_activation_25_16;
wire signed[15:0]    reg_activation_25_17;
wire signed[15:0]    reg_activation_25_18;
wire signed[15:0]    reg_activation_25_19;
wire signed[15:0]    reg_activation_25_20;
wire signed[15:0]    reg_activation_25_21;
wire signed[15:0]    reg_activation_25_22;
wire signed[15:0]    reg_activation_25_23;
wire signed[15:0]    reg_activation_25_24;
wire signed[15:0]    reg_activation_25_25;
wire signed[15:0]    reg_activation_25_26;
wire signed[15:0]    reg_activation_25_27;
wire signed[15:0]    reg_activation_25_28;
wire signed[15:0]    reg_activation_25_29;
wire signed[15:0]    reg_activation_25_30;
wire signed[15:0]    reg_activation_25_31;
wire signed[15:0]    reg_activation_26_0;
wire signed[15:0]    reg_activation_26_1;
wire signed[15:0]    reg_activation_26_2;
wire signed[15:0]    reg_activation_26_3;
wire signed[15:0]    reg_activation_26_4;
wire signed[15:0]    reg_activation_26_5;
wire signed[15:0]    reg_activation_26_6;
wire signed[15:0]    reg_activation_26_7;
wire signed[15:0]    reg_activation_26_8;
wire signed[15:0]    reg_activation_26_9;
wire signed[15:0]    reg_activation_26_10;
wire signed[15:0]    reg_activation_26_11;
wire signed[15:0]    reg_activation_26_12;
wire signed[15:0]    reg_activation_26_13;
wire signed[15:0]    reg_activation_26_14;
wire signed[15:0]    reg_activation_26_15;
wire signed[15:0]    reg_activation_26_16;
wire signed[15:0]    reg_activation_26_17;
wire signed[15:0]    reg_activation_26_18;
wire signed[15:0]    reg_activation_26_19;
wire signed[15:0]    reg_activation_26_20;
wire signed[15:0]    reg_activation_26_21;
wire signed[15:0]    reg_activation_26_22;
wire signed[15:0]    reg_activation_26_23;
wire signed[15:0]    reg_activation_26_24;
wire signed[15:0]    reg_activation_26_25;
wire signed[15:0]    reg_activation_26_26;
wire signed[15:0]    reg_activation_26_27;
wire signed[15:0]    reg_activation_26_28;
wire signed[15:0]    reg_activation_26_29;
wire signed[15:0]    reg_activation_26_30;
wire signed[15:0]    reg_activation_26_31;
wire signed[15:0]    reg_activation_27_0;
wire signed[15:0]    reg_activation_27_1;
wire signed[15:0]    reg_activation_27_2;
wire signed[15:0]    reg_activation_27_3;
wire signed[15:0]    reg_activation_27_4;
wire signed[15:0]    reg_activation_27_5;
wire signed[15:0]    reg_activation_27_6;
wire signed[15:0]    reg_activation_27_7;
wire signed[15:0]    reg_activation_27_8;
wire signed[15:0]    reg_activation_27_9;
wire signed[15:0]    reg_activation_27_10;
wire signed[15:0]    reg_activation_27_11;
wire signed[15:0]    reg_activation_27_12;
wire signed[15:0]    reg_activation_27_13;
wire signed[15:0]    reg_activation_27_14;
wire signed[15:0]    reg_activation_27_15;
wire signed[15:0]    reg_activation_27_16;
wire signed[15:0]    reg_activation_27_17;
wire signed[15:0]    reg_activation_27_18;
wire signed[15:0]    reg_activation_27_19;
wire signed[15:0]    reg_activation_27_20;
wire signed[15:0]    reg_activation_27_21;
wire signed[15:0]    reg_activation_27_22;
wire signed[15:0]    reg_activation_27_23;
wire signed[15:0]    reg_activation_27_24;
wire signed[15:0]    reg_activation_27_25;
wire signed[15:0]    reg_activation_27_26;
wire signed[15:0]    reg_activation_27_27;
wire signed[15:0]    reg_activation_27_28;
wire signed[15:0]    reg_activation_27_29;
wire signed[15:0]    reg_activation_27_30;
wire signed[15:0]    reg_activation_27_31;
wire signed[15:0]    reg_activation_28_0;
wire signed[15:0]    reg_activation_28_1;
wire signed[15:0]    reg_activation_28_2;
wire signed[15:0]    reg_activation_28_3;
wire signed[15:0]    reg_activation_28_4;
wire signed[15:0]    reg_activation_28_5;
wire signed[15:0]    reg_activation_28_6;
wire signed[15:0]    reg_activation_28_7;
wire signed[15:0]    reg_activation_28_8;
wire signed[15:0]    reg_activation_28_9;
wire signed[15:0]    reg_activation_28_10;
wire signed[15:0]    reg_activation_28_11;
wire signed[15:0]    reg_activation_28_12;
wire signed[15:0]    reg_activation_28_13;
wire signed[15:0]    reg_activation_28_14;
wire signed[15:0]    reg_activation_28_15;
wire signed[15:0]    reg_activation_28_16;
wire signed[15:0]    reg_activation_28_17;
wire signed[15:0]    reg_activation_28_18;
wire signed[15:0]    reg_activation_28_19;
wire signed[15:0]    reg_activation_28_20;
wire signed[15:0]    reg_activation_28_21;
wire signed[15:0]    reg_activation_28_22;
wire signed[15:0]    reg_activation_28_23;
wire signed[15:0]    reg_activation_28_24;
wire signed[15:0]    reg_activation_28_25;
wire signed[15:0]    reg_activation_28_26;
wire signed[15:0]    reg_activation_28_27;
wire signed[15:0]    reg_activation_28_28;
wire signed[15:0]    reg_activation_28_29;
wire signed[15:0]    reg_activation_28_30;
wire signed[15:0]    reg_activation_28_31;
wire signed[15:0]    reg_activation_29_0;
wire signed[15:0]    reg_activation_29_1;
wire signed[15:0]    reg_activation_29_2;
wire signed[15:0]    reg_activation_29_3;
wire signed[15:0]    reg_activation_29_4;
wire signed[15:0]    reg_activation_29_5;
wire signed[15:0]    reg_activation_29_6;
wire signed[15:0]    reg_activation_29_7;
wire signed[15:0]    reg_activation_29_8;
wire signed[15:0]    reg_activation_29_9;
wire signed[15:0]    reg_activation_29_10;
wire signed[15:0]    reg_activation_29_11;
wire signed[15:0]    reg_activation_29_12;
wire signed[15:0]    reg_activation_29_13;
wire signed[15:0]    reg_activation_29_14;
wire signed[15:0]    reg_activation_29_15;
wire signed[15:0]    reg_activation_29_16;
wire signed[15:0]    reg_activation_29_17;
wire signed[15:0]    reg_activation_29_18;
wire signed[15:0]    reg_activation_29_19;
wire signed[15:0]    reg_activation_29_20;
wire signed[15:0]    reg_activation_29_21;
wire signed[15:0]    reg_activation_29_22;
wire signed[15:0]    reg_activation_29_23;
wire signed[15:0]    reg_activation_29_24;
wire signed[15:0]    reg_activation_29_25;
wire signed[15:0]    reg_activation_29_26;
wire signed[15:0]    reg_activation_29_27;
wire signed[15:0]    reg_activation_29_28;
wire signed[15:0]    reg_activation_29_29;
wire signed[15:0]    reg_activation_29_30;
wire signed[15:0]    reg_activation_29_31;
wire signed[15:0]    reg_activation_30_0;
wire signed[15:0]    reg_activation_30_1;
wire signed[15:0]    reg_activation_30_2;
wire signed[15:0]    reg_activation_30_3;
wire signed[15:0]    reg_activation_30_4;
wire signed[15:0]    reg_activation_30_5;
wire signed[15:0]    reg_activation_30_6;
wire signed[15:0]    reg_activation_30_7;
wire signed[15:0]    reg_activation_30_8;
wire signed[15:0]    reg_activation_30_9;
wire signed[15:0]    reg_activation_30_10;
wire signed[15:0]    reg_activation_30_11;
wire signed[15:0]    reg_activation_30_12;
wire signed[15:0]    reg_activation_30_13;
wire signed[15:0]    reg_activation_30_14;
wire signed[15:0]    reg_activation_30_15;
wire signed[15:0]    reg_activation_30_16;
wire signed[15:0]    reg_activation_30_17;
wire signed[15:0]    reg_activation_30_18;
wire signed[15:0]    reg_activation_30_19;
wire signed[15:0]    reg_activation_30_20;
wire signed[15:0]    reg_activation_30_21;
wire signed[15:0]    reg_activation_30_22;
wire signed[15:0]    reg_activation_30_23;
wire signed[15:0]    reg_activation_30_24;
wire signed[15:0]    reg_activation_30_25;
wire signed[15:0]    reg_activation_30_26;
wire signed[15:0]    reg_activation_30_27;
wire signed[15:0]    reg_activation_30_28;
wire signed[15:0]    reg_activation_30_29;
wire signed[15:0]    reg_activation_30_30;
wire signed[15:0]    reg_activation_30_31;
wire signed[15:0]    reg_activation_31_0;
wire signed[15:0]    reg_activation_31_1;
wire signed[15:0]    reg_activation_31_2;
wire signed[15:0]    reg_activation_31_3;
wire signed[15:0]    reg_activation_31_4;
wire signed[15:0]    reg_activation_31_5;
wire signed[15:0]    reg_activation_31_6;
wire signed[15:0]    reg_activation_31_7;
wire signed[15:0]    reg_activation_31_8;
wire signed[15:0]    reg_activation_31_9;
wire signed[15:0]    reg_activation_31_10;
wire signed[15:0]    reg_activation_31_11;
wire signed[15:0]    reg_activation_31_12;
wire signed[15:0]    reg_activation_31_13;
wire signed[15:0]    reg_activation_31_14;
wire signed[15:0]    reg_activation_31_15;
wire signed[15:0]    reg_activation_31_16;
wire signed[15:0]    reg_activation_31_17;
wire signed[15:0]    reg_activation_31_18;
wire signed[15:0]    reg_activation_31_19;
wire signed[15:0]    reg_activation_31_20;
wire signed[15:0]    reg_activation_31_21;
wire signed[15:0]    reg_activation_31_22;
wire signed[15:0]    reg_activation_31_23;
wire signed[15:0]    reg_activation_31_24;
wire signed[15:0]    reg_activation_31_25;
wire signed[15:0]    reg_activation_31_26;
wire signed[15:0]    reg_activation_31_27;
wire signed[15:0]    reg_activation_31_28;
wire signed[15:0]    reg_activation_31_29;
wire signed[15:0]    reg_activation_31_30;
wire signed[15:0]    reg_activation_31_31;
wire signed[15:0]    reg_weight_0_0;
wire signed[15:0]    reg_psum_0_0;
wire signed[15:0]    reg_weight_0_1;
wire signed[15:0]    reg_psum_0_1;
wire signed[15:0]    reg_weight_0_2;
wire signed[15:0]    reg_psum_0_2;
wire signed[15:0]    reg_weight_0_3;
wire signed[15:0]    reg_psum_0_3;
wire signed[15:0]    reg_weight_0_4;
wire signed[15:0]    reg_psum_0_4;
wire signed[15:0]    reg_weight_0_5;
wire signed[15:0]    reg_psum_0_5;
wire signed[15:0]    reg_weight_0_6;
wire signed[15:0]    reg_psum_0_6;
wire signed[15:0]    reg_weight_0_7;
wire signed[15:0]    reg_psum_0_7;
wire signed[15:0]    reg_weight_0_8;
wire signed[15:0]    reg_psum_0_8;
wire signed[15:0]    reg_weight_0_9;
wire signed[15:0]    reg_psum_0_9;
wire signed[15:0]    reg_weight_0_10;
wire signed[15:0]    reg_psum_0_10;
wire signed[15:0]    reg_weight_0_11;
wire signed[15:0]    reg_psum_0_11;
wire signed[15:0]    reg_weight_0_12;
wire signed[15:0]    reg_psum_0_12;
wire signed[15:0]    reg_weight_0_13;
wire signed[15:0]    reg_psum_0_13;
wire signed[15:0]    reg_weight_0_14;
wire signed[15:0]    reg_psum_0_14;
wire signed[15:0]    reg_weight_0_15;
wire signed[15:0]    reg_psum_0_15;
wire signed[15:0]    reg_weight_0_16;
wire signed[15:0]    reg_psum_0_16;
wire signed[15:0]    reg_weight_0_17;
wire signed[15:0]    reg_psum_0_17;
wire signed[15:0]    reg_weight_0_18;
wire signed[15:0]    reg_psum_0_18;
wire signed[15:0]    reg_weight_0_19;
wire signed[15:0]    reg_psum_0_19;
wire signed[15:0]    reg_weight_0_20;
wire signed[15:0]    reg_psum_0_20;
wire signed[15:0]    reg_weight_0_21;
wire signed[15:0]    reg_psum_0_21;
wire signed[15:0]    reg_weight_0_22;
wire signed[15:0]    reg_psum_0_22;
wire signed[15:0]    reg_weight_0_23;
wire signed[15:0]    reg_psum_0_23;
wire signed[15:0]    reg_weight_0_24;
wire signed[15:0]    reg_psum_0_24;
wire signed[15:0]    reg_weight_0_25;
wire signed[15:0]    reg_psum_0_25;
wire signed[15:0]    reg_weight_0_26;
wire signed[15:0]    reg_psum_0_26;
wire signed[15:0]    reg_weight_0_27;
wire signed[15:0]    reg_psum_0_27;
wire signed[15:0]    reg_weight_0_28;
wire signed[15:0]    reg_psum_0_28;
wire signed[15:0]    reg_weight_0_29;
wire signed[15:0]    reg_psum_0_29;
wire signed[15:0]    reg_weight_0_30;
wire signed[15:0]    reg_psum_0_30;
wire signed[15:0]    reg_weight_0_31;
wire signed[15:0]    reg_psum_0_31;
wire signed[15:0]    reg_weight_1_0;
wire signed[15:0]    reg_psum_1_0;
wire signed[15:0]    reg_weight_1_1;
wire signed[15:0]    reg_psum_1_1;
wire signed[15:0]    reg_weight_1_2;
wire signed[15:0]    reg_psum_1_2;
wire signed[15:0]    reg_weight_1_3;
wire signed[15:0]    reg_psum_1_3;
wire signed[15:0]    reg_weight_1_4;
wire signed[15:0]    reg_psum_1_4;
wire signed[15:0]    reg_weight_1_5;
wire signed[15:0]    reg_psum_1_5;
wire signed[15:0]    reg_weight_1_6;
wire signed[15:0]    reg_psum_1_6;
wire signed[15:0]    reg_weight_1_7;
wire signed[15:0]    reg_psum_1_7;
wire signed[15:0]    reg_weight_1_8;
wire signed[15:0]    reg_psum_1_8;
wire signed[15:0]    reg_weight_1_9;
wire signed[15:0]    reg_psum_1_9;
wire signed[15:0]    reg_weight_1_10;
wire signed[15:0]    reg_psum_1_10;
wire signed[15:0]    reg_weight_1_11;
wire signed[15:0]    reg_psum_1_11;
wire signed[15:0]    reg_weight_1_12;
wire signed[15:0]    reg_psum_1_12;
wire signed[15:0]    reg_weight_1_13;
wire signed[15:0]    reg_psum_1_13;
wire signed[15:0]    reg_weight_1_14;
wire signed[15:0]    reg_psum_1_14;
wire signed[15:0]    reg_weight_1_15;
wire signed[15:0]    reg_psum_1_15;
wire signed[15:0]    reg_weight_1_16;
wire signed[15:0]    reg_psum_1_16;
wire signed[15:0]    reg_weight_1_17;
wire signed[15:0]    reg_psum_1_17;
wire signed[15:0]    reg_weight_1_18;
wire signed[15:0]    reg_psum_1_18;
wire signed[15:0]    reg_weight_1_19;
wire signed[15:0]    reg_psum_1_19;
wire signed[15:0]    reg_weight_1_20;
wire signed[15:0]    reg_psum_1_20;
wire signed[15:0]    reg_weight_1_21;
wire signed[15:0]    reg_psum_1_21;
wire signed[15:0]    reg_weight_1_22;
wire signed[15:0]    reg_psum_1_22;
wire signed[15:0]    reg_weight_1_23;
wire signed[15:0]    reg_psum_1_23;
wire signed[15:0]    reg_weight_1_24;
wire signed[15:0]    reg_psum_1_24;
wire signed[15:0]    reg_weight_1_25;
wire signed[15:0]    reg_psum_1_25;
wire signed[15:0]    reg_weight_1_26;
wire signed[15:0]    reg_psum_1_26;
wire signed[15:0]    reg_weight_1_27;
wire signed[15:0]    reg_psum_1_27;
wire signed[15:0]    reg_weight_1_28;
wire signed[15:0]    reg_psum_1_28;
wire signed[15:0]    reg_weight_1_29;
wire signed[15:0]    reg_psum_1_29;
wire signed[15:0]    reg_weight_1_30;
wire signed[15:0]    reg_psum_1_30;
wire signed[15:0]    reg_weight_1_31;
wire signed[15:0]    reg_psum_1_31;
wire signed[15:0]    reg_weight_2_0;
wire signed[15:0]    reg_psum_2_0;
wire signed[15:0]    reg_weight_2_1;
wire signed[15:0]    reg_psum_2_1;
wire signed[15:0]    reg_weight_2_2;
wire signed[15:0]    reg_psum_2_2;
wire signed[15:0]    reg_weight_2_3;
wire signed[15:0]    reg_psum_2_3;
wire signed[15:0]    reg_weight_2_4;
wire signed[15:0]    reg_psum_2_4;
wire signed[15:0]    reg_weight_2_5;
wire signed[15:0]    reg_psum_2_5;
wire signed[15:0]    reg_weight_2_6;
wire signed[15:0]    reg_psum_2_6;
wire signed[15:0]    reg_weight_2_7;
wire signed[15:0]    reg_psum_2_7;
wire signed[15:0]    reg_weight_2_8;
wire signed[15:0]    reg_psum_2_8;
wire signed[15:0]    reg_weight_2_9;
wire signed[15:0]    reg_psum_2_9;
wire signed[15:0]    reg_weight_2_10;
wire signed[15:0]    reg_psum_2_10;
wire signed[15:0]    reg_weight_2_11;
wire signed[15:0]    reg_psum_2_11;
wire signed[15:0]    reg_weight_2_12;
wire signed[15:0]    reg_psum_2_12;
wire signed[15:0]    reg_weight_2_13;
wire signed[15:0]    reg_psum_2_13;
wire signed[15:0]    reg_weight_2_14;
wire signed[15:0]    reg_psum_2_14;
wire signed[15:0]    reg_weight_2_15;
wire signed[15:0]    reg_psum_2_15;
wire signed[15:0]    reg_weight_2_16;
wire signed[15:0]    reg_psum_2_16;
wire signed[15:0]    reg_weight_2_17;
wire signed[15:0]    reg_psum_2_17;
wire signed[15:0]    reg_weight_2_18;
wire signed[15:0]    reg_psum_2_18;
wire signed[15:0]    reg_weight_2_19;
wire signed[15:0]    reg_psum_2_19;
wire signed[15:0]    reg_weight_2_20;
wire signed[15:0]    reg_psum_2_20;
wire signed[15:0]    reg_weight_2_21;
wire signed[15:0]    reg_psum_2_21;
wire signed[15:0]    reg_weight_2_22;
wire signed[15:0]    reg_psum_2_22;
wire signed[15:0]    reg_weight_2_23;
wire signed[15:0]    reg_psum_2_23;
wire signed[15:0]    reg_weight_2_24;
wire signed[15:0]    reg_psum_2_24;
wire signed[15:0]    reg_weight_2_25;
wire signed[15:0]    reg_psum_2_25;
wire signed[15:0]    reg_weight_2_26;
wire signed[15:0]    reg_psum_2_26;
wire signed[15:0]    reg_weight_2_27;
wire signed[15:0]    reg_psum_2_27;
wire signed[15:0]    reg_weight_2_28;
wire signed[15:0]    reg_psum_2_28;
wire signed[15:0]    reg_weight_2_29;
wire signed[15:0]    reg_psum_2_29;
wire signed[15:0]    reg_weight_2_30;
wire signed[15:0]    reg_psum_2_30;
wire signed[15:0]    reg_weight_2_31;
wire signed[15:0]    reg_psum_2_31;
wire signed[15:0]    reg_weight_3_0;
wire signed[15:0]    reg_psum_3_0;
wire signed[15:0]    reg_weight_3_1;
wire signed[15:0]    reg_psum_3_1;
wire signed[15:0]    reg_weight_3_2;
wire signed[15:0]    reg_psum_3_2;
wire signed[15:0]    reg_weight_3_3;
wire signed[15:0]    reg_psum_3_3;
wire signed[15:0]    reg_weight_3_4;
wire signed[15:0]    reg_psum_3_4;
wire signed[15:0]    reg_weight_3_5;
wire signed[15:0]    reg_psum_3_5;
wire signed[15:0]    reg_weight_3_6;
wire signed[15:0]    reg_psum_3_6;
wire signed[15:0]    reg_weight_3_7;
wire signed[15:0]    reg_psum_3_7;
wire signed[15:0]    reg_weight_3_8;
wire signed[15:0]    reg_psum_3_8;
wire signed[15:0]    reg_weight_3_9;
wire signed[15:0]    reg_psum_3_9;
wire signed[15:0]    reg_weight_3_10;
wire signed[15:0]    reg_psum_3_10;
wire signed[15:0]    reg_weight_3_11;
wire signed[15:0]    reg_psum_3_11;
wire signed[15:0]    reg_weight_3_12;
wire signed[15:0]    reg_psum_3_12;
wire signed[15:0]    reg_weight_3_13;
wire signed[15:0]    reg_psum_3_13;
wire signed[15:0]    reg_weight_3_14;
wire signed[15:0]    reg_psum_3_14;
wire signed[15:0]    reg_weight_3_15;
wire signed[15:0]    reg_psum_3_15;
wire signed[15:0]    reg_weight_3_16;
wire signed[15:0]    reg_psum_3_16;
wire signed[15:0]    reg_weight_3_17;
wire signed[15:0]    reg_psum_3_17;
wire signed[15:0]    reg_weight_3_18;
wire signed[15:0]    reg_psum_3_18;
wire signed[15:0]    reg_weight_3_19;
wire signed[15:0]    reg_psum_3_19;
wire signed[15:0]    reg_weight_3_20;
wire signed[15:0]    reg_psum_3_20;
wire signed[15:0]    reg_weight_3_21;
wire signed[15:0]    reg_psum_3_21;
wire signed[15:0]    reg_weight_3_22;
wire signed[15:0]    reg_psum_3_22;
wire signed[15:0]    reg_weight_3_23;
wire signed[15:0]    reg_psum_3_23;
wire signed[15:0]    reg_weight_3_24;
wire signed[15:0]    reg_psum_3_24;
wire signed[15:0]    reg_weight_3_25;
wire signed[15:0]    reg_psum_3_25;
wire signed[15:0]    reg_weight_3_26;
wire signed[15:0]    reg_psum_3_26;
wire signed[15:0]    reg_weight_3_27;
wire signed[15:0]    reg_psum_3_27;
wire signed[15:0]    reg_weight_3_28;
wire signed[15:0]    reg_psum_3_28;
wire signed[15:0]    reg_weight_3_29;
wire signed[15:0]    reg_psum_3_29;
wire signed[15:0]    reg_weight_3_30;
wire signed[15:0]    reg_psum_3_30;
wire signed[15:0]    reg_weight_3_31;
wire signed[15:0]    reg_psum_3_31;
wire signed[15:0]    reg_weight_4_0;
wire signed[15:0]    reg_psum_4_0;
wire signed[15:0]    reg_weight_4_1;
wire signed[15:0]    reg_psum_4_1;
wire signed[15:0]    reg_weight_4_2;
wire signed[15:0]    reg_psum_4_2;
wire signed[15:0]    reg_weight_4_3;
wire signed[15:0]    reg_psum_4_3;
wire signed[15:0]    reg_weight_4_4;
wire signed[15:0]    reg_psum_4_4;
wire signed[15:0]    reg_weight_4_5;
wire signed[15:0]    reg_psum_4_5;
wire signed[15:0]    reg_weight_4_6;
wire signed[15:0]    reg_psum_4_6;
wire signed[15:0]    reg_weight_4_7;
wire signed[15:0]    reg_psum_4_7;
wire signed[15:0]    reg_weight_4_8;
wire signed[15:0]    reg_psum_4_8;
wire signed[15:0]    reg_weight_4_9;
wire signed[15:0]    reg_psum_4_9;
wire signed[15:0]    reg_weight_4_10;
wire signed[15:0]    reg_psum_4_10;
wire signed[15:0]    reg_weight_4_11;
wire signed[15:0]    reg_psum_4_11;
wire signed[15:0]    reg_weight_4_12;
wire signed[15:0]    reg_psum_4_12;
wire signed[15:0]    reg_weight_4_13;
wire signed[15:0]    reg_psum_4_13;
wire signed[15:0]    reg_weight_4_14;
wire signed[15:0]    reg_psum_4_14;
wire signed[15:0]    reg_weight_4_15;
wire signed[15:0]    reg_psum_4_15;
wire signed[15:0]    reg_weight_4_16;
wire signed[15:0]    reg_psum_4_16;
wire signed[15:0]    reg_weight_4_17;
wire signed[15:0]    reg_psum_4_17;
wire signed[15:0]    reg_weight_4_18;
wire signed[15:0]    reg_psum_4_18;
wire signed[15:0]    reg_weight_4_19;
wire signed[15:0]    reg_psum_4_19;
wire signed[15:0]    reg_weight_4_20;
wire signed[15:0]    reg_psum_4_20;
wire signed[15:0]    reg_weight_4_21;
wire signed[15:0]    reg_psum_4_21;
wire signed[15:0]    reg_weight_4_22;
wire signed[15:0]    reg_psum_4_22;
wire signed[15:0]    reg_weight_4_23;
wire signed[15:0]    reg_psum_4_23;
wire signed[15:0]    reg_weight_4_24;
wire signed[15:0]    reg_psum_4_24;
wire signed[15:0]    reg_weight_4_25;
wire signed[15:0]    reg_psum_4_25;
wire signed[15:0]    reg_weight_4_26;
wire signed[15:0]    reg_psum_4_26;
wire signed[15:0]    reg_weight_4_27;
wire signed[15:0]    reg_psum_4_27;
wire signed[15:0]    reg_weight_4_28;
wire signed[15:0]    reg_psum_4_28;
wire signed[15:0]    reg_weight_4_29;
wire signed[15:0]    reg_psum_4_29;
wire signed[15:0]    reg_weight_4_30;
wire signed[15:0]    reg_psum_4_30;
wire signed[15:0]    reg_weight_4_31;
wire signed[15:0]    reg_psum_4_31;
wire signed[15:0]    reg_weight_5_0;
wire signed[15:0]    reg_psum_5_0;
wire signed[15:0]    reg_weight_5_1;
wire signed[15:0]    reg_psum_5_1;
wire signed[15:0]    reg_weight_5_2;
wire signed[15:0]    reg_psum_5_2;
wire signed[15:0]    reg_weight_5_3;
wire signed[15:0]    reg_psum_5_3;
wire signed[15:0]    reg_weight_5_4;
wire signed[15:0]    reg_psum_5_4;
wire signed[15:0]    reg_weight_5_5;
wire signed[15:0]    reg_psum_5_5;
wire signed[15:0]    reg_weight_5_6;
wire signed[15:0]    reg_psum_5_6;
wire signed[15:0]    reg_weight_5_7;
wire signed[15:0]    reg_psum_5_7;
wire signed[15:0]    reg_weight_5_8;
wire signed[15:0]    reg_psum_5_8;
wire signed[15:0]    reg_weight_5_9;
wire signed[15:0]    reg_psum_5_9;
wire signed[15:0]    reg_weight_5_10;
wire signed[15:0]    reg_psum_5_10;
wire signed[15:0]    reg_weight_5_11;
wire signed[15:0]    reg_psum_5_11;
wire signed[15:0]    reg_weight_5_12;
wire signed[15:0]    reg_psum_5_12;
wire signed[15:0]    reg_weight_5_13;
wire signed[15:0]    reg_psum_5_13;
wire signed[15:0]    reg_weight_5_14;
wire signed[15:0]    reg_psum_5_14;
wire signed[15:0]    reg_weight_5_15;
wire signed[15:0]    reg_psum_5_15;
wire signed[15:0]    reg_weight_5_16;
wire signed[15:0]    reg_psum_5_16;
wire signed[15:0]    reg_weight_5_17;
wire signed[15:0]    reg_psum_5_17;
wire signed[15:0]    reg_weight_5_18;
wire signed[15:0]    reg_psum_5_18;
wire signed[15:0]    reg_weight_5_19;
wire signed[15:0]    reg_psum_5_19;
wire signed[15:0]    reg_weight_5_20;
wire signed[15:0]    reg_psum_5_20;
wire signed[15:0]    reg_weight_5_21;
wire signed[15:0]    reg_psum_5_21;
wire signed[15:0]    reg_weight_5_22;
wire signed[15:0]    reg_psum_5_22;
wire signed[15:0]    reg_weight_5_23;
wire signed[15:0]    reg_psum_5_23;
wire signed[15:0]    reg_weight_5_24;
wire signed[15:0]    reg_psum_5_24;
wire signed[15:0]    reg_weight_5_25;
wire signed[15:0]    reg_psum_5_25;
wire signed[15:0]    reg_weight_5_26;
wire signed[15:0]    reg_psum_5_26;
wire signed[15:0]    reg_weight_5_27;
wire signed[15:0]    reg_psum_5_27;
wire signed[15:0]    reg_weight_5_28;
wire signed[15:0]    reg_psum_5_28;
wire signed[15:0]    reg_weight_5_29;
wire signed[15:0]    reg_psum_5_29;
wire signed[15:0]    reg_weight_5_30;
wire signed[15:0]    reg_psum_5_30;
wire signed[15:0]    reg_weight_5_31;
wire signed[15:0]    reg_psum_5_31;
wire signed[15:0]    reg_weight_6_0;
wire signed[15:0]    reg_psum_6_0;
wire signed[15:0]    reg_weight_6_1;
wire signed[15:0]    reg_psum_6_1;
wire signed[15:0]    reg_weight_6_2;
wire signed[15:0]    reg_psum_6_2;
wire signed[15:0]    reg_weight_6_3;
wire signed[15:0]    reg_psum_6_3;
wire signed[15:0]    reg_weight_6_4;
wire signed[15:0]    reg_psum_6_4;
wire signed[15:0]    reg_weight_6_5;
wire signed[15:0]    reg_psum_6_5;
wire signed[15:0]    reg_weight_6_6;
wire signed[15:0]    reg_psum_6_6;
wire signed[15:0]    reg_weight_6_7;
wire signed[15:0]    reg_psum_6_7;
wire signed[15:0]    reg_weight_6_8;
wire signed[15:0]    reg_psum_6_8;
wire signed[15:0]    reg_weight_6_9;
wire signed[15:0]    reg_psum_6_9;
wire signed[15:0]    reg_weight_6_10;
wire signed[15:0]    reg_psum_6_10;
wire signed[15:0]    reg_weight_6_11;
wire signed[15:0]    reg_psum_6_11;
wire signed[15:0]    reg_weight_6_12;
wire signed[15:0]    reg_psum_6_12;
wire signed[15:0]    reg_weight_6_13;
wire signed[15:0]    reg_psum_6_13;
wire signed[15:0]    reg_weight_6_14;
wire signed[15:0]    reg_psum_6_14;
wire signed[15:0]    reg_weight_6_15;
wire signed[15:0]    reg_psum_6_15;
wire signed[15:0]    reg_weight_6_16;
wire signed[15:0]    reg_psum_6_16;
wire signed[15:0]    reg_weight_6_17;
wire signed[15:0]    reg_psum_6_17;
wire signed[15:0]    reg_weight_6_18;
wire signed[15:0]    reg_psum_6_18;
wire signed[15:0]    reg_weight_6_19;
wire signed[15:0]    reg_psum_6_19;
wire signed[15:0]    reg_weight_6_20;
wire signed[15:0]    reg_psum_6_20;
wire signed[15:0]    reg_weight_6_21;
wire signed[15:0]    reg_psum_6_21;
wire signed[15:0]    reg_weight_6_22;
wire signed[15:0]    reg_psum_6_22;
wire signed[15:0]    reg_weight_6_23;
wire signed[15:0]    reg_psum_6_23;
wire signed[15:0]    reg_weight_6_24;
wire signed[15:0]    reg_psum_6_24;
wire signed[15:0]    reg_weight_6_25;
wire signed[15:0]    reg_psum_6_25;
wire signed[15:0]    reg_weight_6_26;
wire signed[15:0]    reg_psum_6_26;
wire signed[15:0]    reg_weight_6_27;
wire signed[15:0]    reg_psum_6_27;
wire signed[15:0]    reg_weight_6_28;
wire signed[15:0]    reg_psum_6_28;
wire signed[15:0]    reg_weight_6_29;
wire signed[15:0]    reg_psum_6_29;
wire signed[15:0]    reg_weight_6_30;
wire signed[15:0]    reg_psum_6_30;
wire signed[15:0]    reg_weight_6_31;
wire signed[15:0]    reg_psum_6_31;
wire signed[15:0]    reg_weight_7_0;
wire signed[15:0]    reg_psum_7_0;
wire signed[15:0]    reg_weight_7_1;
wire signed[15:0]    reg_psum_7_1;
wire signed[15:0]    reg_weight_7_2;
wire signed[15:0]    reg_psum_7_2;
wire signed[15:0]    reg_weight_7_3;
wire signed[15:0]    reg_psum_7_3;
wire signed[15:0]    reg_weight_7_4;
wire signed[15:0]    reg_psum_7_4;
wire signed[15:0]    reg_weight_7_5;
wire signed[15:0]    reg_psum_7_5;
wire signed[15:0]    reg_weight_7_6;
wire signed[15:0]    reg_psum_7_6;
wire signed[15:0]    reg_weight_7_7;
wire signed[15:0]    reg_psum_7_7;
wire signed[15:0]    reg_weight_7_8;
wire signed[15:0]    reg_psum_7_8;
wire signed[15:0]    reg_weight_7_9;
wire signed[15:0]    reg_psum_7_9;
wire signed[15:0]    reg_weight_7_10;
wire signed[15:0]    reg_psum_7_10;
wire signed[15:0]    reg_weight_7_11;
wire signed[15:0]    reg_psum_7_11;
wire signed[15:0]    reg_weight_7_12;
wire signed[15:0]    reg_psum_7_12;
wire signed[15:0]    reg_weight_7_13;
wire signed[15:0]    reg_psum_7_13;
wire signed[15:0]    reg_weight_7_14;
wire signed[15:0]    reg_psum_7_14;
wire signed[15:0]    reg_weight_7_15;
wire signed[15:0]    reg_psum_7_15;
wire signed[15:0]    reg_weight_7_16;
wire signed[15:0]    reg_psum_7_16;
wire signed[15:0]    reg_weight_7_17;
wire signed[15:0]    reg_psum_7_17;
wire signed[15:0]    reg_weight_7_18;
wire signed[15:0]    reg_psum_7_18;
wire signed[15:0]    reg_weight_7_19;
wire signed[15:0]    reg_psum_7_19;
wire signed[15:0]    reg_weight_7_20;
wire signed[15:0]    reg_psum_7_20;
wire signed[15:0]    reg_weight_7_21;
wire signed[15:0]    reg_psum_7_21;
wire signed[15:0]    reg_weight_7_22;
wire signed[15:0]    reg_psum_7_22;
wire signed[15:0]    reg_weight_7_23;
wire signed[15:0]    reg_psum_7_23;
wire signed[15:0]    reg_weight_7_24;
wire signed[15:0]    reg_psum_7_24;
wire signed[15:0]    reg_weight_7_25;
wire signed[15:0]    reg_psum_7_25;
wire signed[15:0]    reg_weight_7_26;
wire signed[15:0]    reg_psum_7_26;
wire signed[15:0]    reg_weight_7_27;
wire signed[15:0]    reg_psum_7_27;
wire signed[15:0]    reg_weight_7_28;
wire signed[15:0]    reg_psum_7_28;
wire signed[15:0]    reg_weight_7_29;
wire signed[15:0]    reg_psum_7_29;
wire signed[15:0]    reg_weight_7_30;
wire signed[15:0]    reg_psum_7_30;
wire signed[15:0]    reg_weight_7_31;
wire signed[15:0]    reg_psum_7_31;
wire signed[15:0]    reg_weight_8_0;
wire signed[15:0]    reg_psum_8_0;
wire signed[15:0]    reg_weight_8_1;
wire signed[15:0]    reg_psum_8_1;
wire signed[15:0]    reg_weight_8_2;
wire signed[15:0]    reg_psum_8_2;
wire signed[15:0]    reg_weight_8_3;
wire signed[15:0]    reg_psum_8_3;
wire signed[15:0]    reg_weight_8_4;
wire signed[15:0]    reg_psum_8_4;
wire signed[15:0]    reg_weight_8_5;
wire signed[15:0]    reg_psum_8_5;
wire signed[15:0]    reg_weight_8_6;
wire signed[15:0]    reg_psum_8_6;
wire signed[15:0]    reg_weight_8_7;
wire signed[15:0]    reg_psum_8_7;
wire signed[15:0]    reg_weight_8_8;
wire signed[15:0]    reg_psum_8_8;
wire signed[15:0]    reg_weight_8_9;
wire signed[15:0]    reg_psum_8_9;
wire signed[15:0]    reg_weight_8_10;
wire signed[15:0]    reg_psum_8_10;
wire signed[15:0]    reg_weight_8_11;
wire signed[15:0]    reg_psum_8_11;
wire signed[15:0]    reg_weight_8_12;
wire signed[15:0]    reg_psum_8_12;
wire signed[15:0]    reg_weight_8_13;
wire signed[15:0]    reg_psum_8_13;
wire signed[15:0]    reg_weight_8_14;
wire signed[15:0]    reg_psum_8_14;
wire signed[15:0]    reg_weight_8_15;
wire signed[15:0]    reg_psum_8_15;
wire signed[15:0]    reg_weight_8_16;
wire signed[15:0]    reg_psum_8_16;
wire signed[15:0]    reg_weight_8_17;
wire signed[15:0]    reg_psum_8_17;
wire signed[15:0]    reg_weight_8_18;
wire signed[15:0]    reg_psum_8_18;
wire signed[15:0]    reg_weight_8_19;
wire signed[15:0]    reg_psum_8_19;
wire signed[15:0]    reg_weight_8_20;
wire signed[15:0]    reg_psum_8_20;
wire signed[15:0]    reg_weight_8_21;
wire signed[15:0]    reg_psum_8_21;
wire signed[15:0]    reg_weight_8_22;
wire signed[15:0]    reg_psum_8_22;
wire signed[15:0]    reg_weight_8_23;
wire signed[15:0]    reg_psum_8_23;
wire signed[15:0]    reg_weight_8_24;
wire signed[15:0]    reg_psum_8_24;
wire signed[15:0]    reg_weight_8_25;
wire signed[15:0]    reg_psum_8_25;
wire signed[15:0]    reg_weight_8_26;
wire signed[15:0]    reg_psum_8_26;
wire signed[15:0]    reg_weight_8_27;
wire signed[15:0]    reg_psum_8_27;
wire signed[15:0]    reg_weight_8_28;
wire signed[15:0]    reg_psum_8_28;
wire signed[15:0]    reg_weight_8_29;
wire signed[15:0]    reg_psum_8_29;
wire signed[15:0]    reg_weight_8_30;
wire signed[15:0]    reg_psum_8_30;
wire signed[15:0]    reg_weight_8_31;
wire signed[15:0]    reg_psum_8_31;
wire signed[15:0]    reg_weight_9_0;
wire signed[15:0]    reg_psum_9_0;
wire signed[15:0]    reg_weight_9_1;
wire signed[15:0]    reg_psum_9_1;
wire signed[15:0]    reg_weight_9_2;
wire signed[15:0]    reg_psum_9_2;
wire signed[15:0]    reg_weight_9_3;
wire signed[15:0]    reg_psum_9_3;
wire signed[15:0]    reg_weight_9_4;
wire signed[15:0]    reg_psum_9_4;
wire signed[15:0]    reg_weight_9_5;
wire signed[15:0]    reg_psum_9_5;
wire signed[15:0]    reg_weight_9_6;
wire signed[15:0]    reg_psum_9_6;
wire signed[15:0]    reg_weight_9_7;
wire signed[15:0]    reg_psum_9_7;
wire signed[15:0]    reg_weight_9_8;
wire signed[15:0]    reg_psum_9_8;
wire signed[15:0]    reg_weight_9_9;
wire signed[15:0]    reg_psum_9_9;
wire signed[15:0]    reg_weight_9_10;
wire signed[15:0]    reg_psum_9_10;
wire signed[15:0]    reg_weight_9_11;
wire signed[15:0]    reg_psum_9_11;
wire signed[15:0]    reg_weight_9_12;
wire signed[15:0]    reg_psum_9_12;
wire signed[15:0]    reg_weight_9_13;
wire signed[15:0]    reg_psum_9_13;
wire signed[15:0]    reg_weight_9_14;
wire signed[15:0]    reg_psum_9_14;
wire signed[15:0]    reg_weight_9_15;
wire signed[15:0]    reg_psum_9_15;
wire signed[15:0]    reg_weight_9_16;
wire signed[15:0]    reg_psum_9_16;
wire signed[15:0]    reg_weight_9_17;
wire signed[15:0]    reg_psum_9_17;
wire signed[15:0]    reg_weight_9_18;
wire signed[15:0]    reg_psum_9_18;
wire signed[15:0]    reg_weight_9_19;
wire signed[15:0]    reg_psum_9_19;
wire signed[15:0]    reg_weight_9_20;
wire signed[15:0]    reg_psum_9_20;
wire signed[15:0]    reg_weight_9_21;
wire signed[15:0]    reg_psum_9_21;
wire signed[15:0]    reg_weight_9_22;
wire signed[15:0]    reg_psum_9_22;
wire signed[15:0]    reg_weight_9_23;
wire signed[15:0]    reg_psum_9_23;
wire signed[15:0]    reg_weight_9_24;
wire signed[15:0]    reg_psum_9_24;
wire signed[15:0]    reg_weight_9_25;
wire signed[15:0]    reg_psum_9_25;
wire signed[15:0]    reg_weight_9_26;
wire signed[15:0]    reg_psum_9_26;
wire signed[15:0]    reg_weight_9_27;
wire signed[15:0]    reg_psum_9_27;
wire signed[15:0]    reg_weight_9_28;
wire signed[15:0]    reg_psum_9_28;
wire signed[15:0]    reg_weight_9_29;
wire signed[15:0]    reg_psum_9_29;
wire signed[15:0]    reg_weight_9_30;
wire signed[15:0]    reg_psum_9_30;
wire signed[15:0]    reg_weight_9_31;
wire signed[15:0]    reg_psum_9_31;
wire signed[15:0]    reg_weight_10_0;
wire signed[15:0]    reg_psum_10_0;
wire signed[15:0]    reg_weight_10_1;
wire signed[15:0]    reg_psum_10_1;
wire signed[15:0]    reg_weight_10_2;
wire signed[15:0]    reg_psum_10_2;
wire signed[15:0]    reg_weight_10_3;
wire signed[15:0]    reg_psum_10_3;
wire signed[15:0]    reg_weight_10_4;
wire signed[15:0]    reg_psum_10_4;
wire signed[15:0]    reg_weight_10_5;
wire signed[15:0]    reg_psum_10_5;
wire signed[15:0]    reg_weight_10_6;
wire signed[15:0]    reg_psum_10_6;
wire signed[15:0]    reg_weight_10_7;
wire signed[15:0]    reg_psum_10_7;
wire signed[15:0]    reg_weight_10_8;
wire signed[15:0]    reg_psum_10_8;
wire signed[15:0]    reg_weight_10_9;
wire signed[15:0]    reg_psum_10_9;
wire signed[15:0]    reg_weight_10_10;
wire signed[15:0]    reg_psum_10_10;
wire signed[15:0]    reg_weight_10_11;
wire signed[15:0]    reg_psum_10_11;
wire signed[15:0]    reg_weight_10_12;
wire signed[15:0]    reg_psum_10_12;
wire signed[15:0]    reg_weight_10_13;
wire signed[15:0]    reg_psum_10_13;
wire signed[15:0]    reg_weight_10_14;
wire signed[15:0]    reg_psum_10_14;
wire signed[15:0]    reg_weight_10_15;
wire signed[15:0]    reg_psum_10_15;
wire signed[15:0]    reg_weight_10_16;
wire signed[15:0]    reg_psum_10_16;
wire signed[15:0]    reg_weight_10_17;
wire signed[15:0]    reg_psum_10_17;
wire signed[15:0]    reg_weight_10_18;
wire signed[15:0]    reg_psum_10_18;
wire signed[15:0]    reg_weight_10_19;
wire signed[15:0]    reg_psum_10_19;
wire signed[15:0]    reg_weight_10_20;
wire signed[15:0]    reg_psum_10_20;
wire signed[15:0]    reg_weight_10_21;
wire signed[15:0]    reg_psum_10_21;
wire signed[15:0]    reg_weight_10_22;
wire signed[15:0]    reg_psum_10_22;
wire signed[15:0]    reg_weight_10_23;
wire signed[15:0]    reg_psum_10_23;
wire signed[15:0]    reg_weight_10_24;
wire signed[15:0]    reg_psum_10_24;
wire signed[15:0]    reg_weight_10_25;
wire signed[15:0]    reg_psum_10_25;
wire signed[15:0]    reg_weight_10_26;
wire signed[15:0]    reg_psum_10_26;
wire signed[15:0]    reg_weight_10_27;
wire signed[15:0]    reg_psum_10_27;
wire signed[15:0]    reg_weight_10_28;
wire signed[15:0]    reg_psum_10_28;
wire signed[15:0]    reg_weight_10_29;
wire signed[15:0]    reg_psum_10_29;
wire signed[15:0]    reg_weight_10_30;
wire signed[15:0]    reg_psum_10_30;
wire signed[15:0]    reg_weight_10_31;
wire signed[15:0]    reg_psum_10_31;
wire signed[15:0]    reg_weight_11_0;
wire signed[15:0]    reg_psum_11_0;
wire signed[15:0]    reg_weight_11_1;
wire signed[15:0]    reg_psum_11_1;
wire signed[15:0]    reg_weight_11_2;
wire signed[15:0]    reg_psum_11_2;
wire signed[15:0]    reg_weight_11_3;
wire signed[15:0]    reg_psum_11_3;
wire signed[15:0]    reg_weight_11_4;
wire signed[15:0]    reg_psum_11_4;
wire signed[15:0]    reg_weight_11_5;
wire signed[15:0]    reg_psum_11_5;
wire signed[15:0]    reg_weight_11_6;
wire signed[15:0]    reg_psum_11_6;
wire signed[15:0]    reg_weight_11_7;
wire signed[15:0]    reg_psum_11_7;
wire signed[15:0]    reg_weight_11_8;
wire signed[15:0]    reg_psum_11_8;
wire signed[15:0]    reg_weight_11_9;
wire signed[15:0]    reg_psum_11_9;
wire signed[15:0]    reg_weight_11_10;
wire signed[15:0]    reg_psum_11_10;
wire signed[15:0]    reg_weight_11_11;
wire signed[15:0]    reg_psum_11_11;
wire signed[15:0]    reg_weight_11_12;
wire signed[15:0]    reg_psum_11_12;
wire signed[15:0]    reg_weight_11_13;
wire signed[15:0]    reg_psum_11_13;
wire signed[15:0]    reg_weight_11_14;
wire signed[15:0]    reg_psum_11_14;
wire signed[15:0]    reg_weight_11_15;
wire signed[15:0]    reg_psum_11_15;
wire signed[15:0]    reg_weight_11_16;
wire signed[15:0]    reg_psum_11_16;
wire signed[15:0]    reg_weight_11_17;
wire signed[15:0]    reg_psum_11_17;
wire signed[15:0]    reg_weight_11_18;
wire signed[15:0]    reg_psum_11_18;
wire signed[15:0]    reg_weight_11_19;
wire signed[15:0]    reg_psum_11_19;
wire signed[15:0]    reg_weight_11_20;
wire signed[15:0]    reg_psum_11_20;
wire signed[15:0]    reg_weight_11_21;
wire signed[15:0]    reg_psum_11_21;
wire signed[15:0]    reg_weight_11_22;
wire signed[15:0]    reg_psum_11_22;
wire signed[15:0]    reg_weight_11_23;
wire signed[15:0]    reg_psum_11_23;
wire signed[15:0]    reg_weight_11_24;
wire signed[15:0]    reg_psum_11_24;
wire signed[15:0]    reg_weight_11_25;
wire signed[15:0]    reg_psum_11_25;
wire signed[15:0]    reg_weight_11_26;
wire signed[15:0]    reg_psum_11_26;
wire signed[15:0]    reg_weight_11_27;
wire signed[15:0]    reg_psum_11_27;
wire signed[15:0]    reg_weight_11_28;
wire signed[15:0]    reg_psum_11_28;
wire signed[15:0]    reg_weight_11_29;
wire signed[15:0]    reg_psum_11_29;
wire signed[15:0]    reg_weight_11_30;
wire signed[15:0]    reg_psum_11_30;
wire signed[15:0]    reg_weight_11_31;
wire signed[15:0]    reg_psum_11_31;
wire signed[15:0]    reg_weight_12_0;
wire signed[15:0]    reg_psum_12_0;
wire signed[15:0]    reg_weight_12_1;
wire signed[15:0]    reg_psum_12_1;
wire signed[15:0]    reg_weight_12_2;
wire signed[15:0]    reg_psum_12_2;
wire signed[15:0]    reg_weight_12_3;
wire signed[15:0]    reg_psum_12_3;
wire signed[15:0]    reg_weight_12_4;
wire signed[15:0]    reg_psum_12_4;
wire signed[15:0]    reg_weight_12_5;
wire signed[15:0]    reg_psum_12_5;
wire signed[15:0]    reg_weight_12_6;
wire signed[15:0]    reg_psum_12_6;
wire signed[15:0]    reg_weight_12_7;
wire signed[15:0]    reg_psum_12_7;
wire signed[15:0]    reg_weight_12_8;
wire signed[15:0]    reg_psum_12_8;
wire signed[15:0]    reg_weight_12_9;
wire signed[15:0]    reg_psum_12_9;
wire signed[15:0]    reg_weight_12_10;
wire signed[15:0]    reg_psum_12_10;
wire signed[15:0]    reg_weight_12_11;
wire signed[15:0]    reg_psum_12_11;
wire signed[15:0]    reg_weight_12_12;
wire signed[15:0]    reg_psum_12_12;
wire signed[15:0]    reg_weight_12_13;
wire signed[15:0]    reg_psum_12_13;
wire signed[15:0]    reg_weight_12_14;
wire signed[15:0]    reg_psum_12_14;
wire signed[15:0]    reg_weight_12_15;
wire signed[15:0]    reg_psum_12_15;
wire signed[15:0]    reg_weight_12_16;
wire signed[15:0]    reg_psum_12_16;
wire signed[15:0]    reg_weight_12_17;
wire signed[15:0]    reg_psum_12_17;
wire signed[15:0]    reg_weight_12_18;
wire signed[15:0]    reg_psum_12_18;
wire signed[15:0]    reg_weight_12_19;
wire signed[15:0]    reg_psum_12_19;
wire signed[15:0]    reg_weight_12_20;
wire signed[15:0]    reg_psum_12_20;
wire signed[15:0]    reg_weight_12_21;
wire signed[15:0]    reg_psum_12_21;
wire signed[15:0]    reg_weight_12_22;
wire signed[15:0]    reg_psum_12_22;
wire signed[15:0]    reg_weight_12_23;
wire signed[15:0]    reg_psum_12_23;
wire signed[15:0]    reg_weight_12_24;
wire signed[15:0]    reg_psum_12_24;
wire signed[15:0]    reg_weight_12_25;
wire signed[15:0]    reg_psum_12_25;
wire signed[15:0]    reg_weight_12_26;
wire signed[15:0]    reg_psum_12_26;
wire signed[15:0]    reg_weight_12_27;
wire signed[15:0]    reg_psum_12_27;
wire signed[15:0]    reg_weight_12_28;
wire signed[15:0]    reg_psum_12_28;
wire signed[15:0]    reg_weight_12_29;
wire signed[15:0]    reg_psum_12_29;
wire signed[15:0]    reg_weight_12_30;
wire signed[15:0]    reg_psum_12_30;
wire signed[15:0]    reg_weight_12_31;
wire signed[15:0]    reg_psum_12_31;
wire signed[15:0]    reg_weight_13_0;
wire signed[15:0]    reg_psum_13_0;
wire signed[15:0]    reg_weight_13_1;
wire signed[15:0]    reg_psum_13_1;
wire signed[15:0]    reg_weight_13_2;
wire signed[15:0]    reg_psum_13_2;
wire signed[15:0]    reg_weight_13_3;
wire signed[15:0]    reg_psum_13_3;
wire signed[15:0]    reg_weight_13_4;
wire signed[15:0]    reg_psum_13_4;
wire signed[15:0]    reg_weight_13_5;
wire signed[15:0]    reg_psum_13_5;
wire signed[15:0]    reg_weight_13_6;
wire signed[15:0]    reg_psum_13_6;
wire signed[15:0]    reg_weight_13_7;
wire signed[15:0]    reg_psum_13_7;
wire signed[15:0]    reg_weight_13_8;
wire signed[15:0]    reg_psum_13_8;
wire signed[15:0]    reg_weight_13_9;
wire signed[15:0]    reg_psum_13_9;
wire signed[15:0]    reg_weight_13_10;
wire signed[15:0]    reg_psum_13_10;
wire signed[15:0]    reg_weight_13_11;
wire signed[15:0]    reg_psum_13_11;
wire signed[15:0]    reg_weight_13_12;
wire signed[15:0]    reg_psum_13_12;
wire signed[15:0]    reg_weight_13_13;
wire signed[15:0]    reg_psum_13_13;
wire signed[15:0]    reg_weight_13_14;
wire signed[15:0]    reg_psum_13_14;
wire signed[15:0]    reg_weight_13_15;
wire signed[15:0]    reg_psum_13_15;
wire signed[15:0]    reg_weight_13_16;
wire signed[15:0]    reg_psum_13_16;
wire signed[15:0]    reg_weight_13_17;
wire signed[15:0]    reg_psum_13_17;
wire signed[15:0]    reg_weight_13_18;
wire signed[15:0]    reg_psum_13_18;
wire signed[15:0]    reg_weight_13_19;
wire signed[15:0]    reg_psum_13_19;
wire signed[15:0]    reg_weight_13_20;
wire signed[15:0]    reg_psum_13_20;
wire signed[15:0]    reg_weight_13_21;
wire signed[15:0]    reg_psum_13_21;
wire signed[15:0]    reg_weight_13_22;
wire signed[15:0]    reg_psum_13_22;
wire signed[15:0]    reg_weight_13_23;
wire signed[15:0]    reg_psum_13_23;
wire signed[15:0]    reg_weight_13_24;
wire signed[15:0]    reg_psum_13_24;
wire signed[15:0]    reg_weight_13_25;
wire signed[15:0]    reg_psum_13_25;
wire signed[15:0]    reg_weight_13_26;
wire signed[15:0]    reg_psum_13_26;
wire signed[15:0]    reg_weight_13_27;
wire signed[15:0]    reg_psum_13_27;
wire signed[15:0]    reg_weight_13_28;
wire signed[15:0]    reg_psum_13_28;
wire signed[15:0]    reg_weight_13_29;
wire signed[15:0]    reg_psum_13_29;
wire signed[15:0]    reg_weight_13_30;
wire signed[15:0]    reg_psum_13_30;
wire signed[15:0]    reg_weight_13_31;
wire signed[15:0]    reg_psum_13_31;
wire signed[15:0]    reg_weight_14_0;
wire signed[15:0]    reg_psum_14_0;
wire signed[15:0]    reg_weight_14_1;
wire signed[15:0]    reg_psum_14_1;
wire signed[15:0]    reg_weight_14_2;
wire signed[15:0]    reg_psum_14_2;
wire signed[15:0]    reg_weight_14_3;
wire signed[15:0]    reg_psum_14_3;
wire signed[15:0]    reg_weight_14_4;
wire signed[15:0]    reg_psum_14_4;
wire signed[15:0]    reg_weight_14_5;
wire signed[15:0]    reg_psum_14_5;
wire signed[15:0]    reg_weight_14_6;
wire signed[15:0]    reg_psum_14_6;
wire signed[15:0]    reg_weight_14_7;
wire signed[15:0]    reg_psum_14_7;
wire signed[15:0]    reg_weight_14_8;
wire signed[15:0]    reg_psum_14_8;
wire signed[15:0]    reg_weight_14_9;
wire signed[15:0]    reg_psum_14_9;
wire signed[15:0]    reg_weight_14_10;
wire signed[15:0]    reg_psum_14_10;
wire signed[15:0]    reg_weight_14_11;
wire signed[15:0]    reg_psum_14_11;
wire signed[15:0]    reg_weight_14_12;
wire signed[15:0]    reg_psum_14_12;
wire signed[15:0]    reg_weight_14_13;
wire signed[15:0]    reg_psum_14_13;
wire signed[15:0]    reg_weight_14_14;
wire signed[15:0]    reg_psum_14_14;
wire signed[15:0]    reg_weight_14_15;
wire signed[15:0]    reg_psum_14_15;
wire signed[15:0]    reg_weight_14_16;
wire signed[15:0]    reg_psum_14_16;
wire signed[15:0]    reg_weight_14_17;
wire signed[15:0]    reg_psum_14_17;
wire signed[15:0]    reg_weight_14_18;
wire signed[15:0]    reg_psum_14_18;
wire signed[15:0]    reg_weight_14_19;
wire signed[15:0]    reg_psum_14_19;
wire signed[15:0]    reg_weight_14_20;
wire signed[15:0]    reg_psum_14_20;
wire signed[15:0]    reg_weight_14_21;
wire signed[15:0]    reg_psum_14_21;
wire signed[15:0]    reg_weight_14_22;
wire signed[15:0]    reg_psum_14_22;
wire signed[15:0]    reg_weight_14_23;
wire signed[15:0]    reg_psum_14_23;
wire signed[15:0]    reg_weight_14_24;
wire signed[15:0]    reg_psum_14_24;
wire signed[15:0]    reg_weight_14_25;
wire signed[15:0]    reg_psum_14_25;
wire signed[15:0]    reg_weight_14_26;
wire signed[15:0]    reg_psum_14_26;
wire signed[15:0]    reg_weight_14_27;
wire signed[15:0]    reg_psum_14_27;
wire signed[15:0]    reg_weight_14_28;
wire signed[15:0]    reg_psum_14_28;
wire signed[15:0]    reg_weight_14_29;
wire signed[15:0]    reg_psum_14_29;
wire signed[15:0]    reg_weight_14_30;
wire signed[15:0]    reg_psum_14_30;
wire signed[15:0]    reg_weight_14_31;
wire signed[15:0]    reg_psum_14_31;
wire signed[15:0]    reg_weight_15_0;
wire signed[15:0]    reg_psum_15_0;
wire signed[15:0]    reg_weight_15_1;
wire signed[15:0]    reg_psum_15_1;
wire signed[15:0]    reg_weight_15_2;
wire signed[15:0]    reg_psum_15_2;
wire signed[15:0]    reg_weight_15_3;
wire signed[15:0]    reg_psum_15_3;
wire signed[15:0]    reg_weight_15_4;
wire signed[15:0]    reg_psum_15_4;
wire signed[15:0]    reg_weight_15_5;
wire signed[15:0]    reg_psum_15_5;
wire signed[15:0]    reg_weight_15_6;
wire signed[15:0]    reg_psum_15_6;
wire signed[15:0]    reg_weight_15_7;
wire signed[15:0]    reg_psum_15_7;
wire signed[15:0]    reg_weight_15_8;
wire signed[15:0]    reg_psum_15_8;
wire signed[15:0]    reg_weight_15_9;
wire signed[15:0]    reg_psum_15_9;
wire signed[15:0]    reg_weight_15_10;
wire signed[15:0]    reg_psum_15_10;
wire signed[15:0]    reg_weight_15_11;
wire signed[15:0]    reg_psum_15_11;
wire signed[15:0]    reg_weight_15_12;
wire signed[15:0]    reg_psum_15_12;
wire signed[15:0]    reg_weight_15_13;
wire signed[15:0]    reg_psum_15_13;
wire signed[15:0]    reg_weight_15_14;
wire signed[15:0]    reg_psum_15_14;
wire signed[15:0]    reg_weight_15_15;
wire signed[15:0]    reg_psum_15_15;
wire signed[15:0]    reg_weight_15_16;
wire signed[15:0]    reg_psum_15_16;
wire signed[15:0]    reg_weight_15_17;
wire signed[15:0]    reg_psum_15_17;
wire signed[15:0]    reg_weight_15_18;
wire signed[15:0]    reg_psum_15_18;
wire signed[15:0]    reg_weight_15_19;
wire signed[15:0]    reg_psum_15_19;
wire signed[15:0]    reg_weight_15_20;
wire signed[15:0]    reg_psum_15_20;
wire signed[15:0]    reg_weight_15_21;
wire signed[15:0]    reg_psum_15_21;
wire signed[15:0]    reg_weight_15_22;
wire signed[15:0]    reg_psum_15_22;
wire signed[15:0]    reg_weight_15_23;
wire signed[15:0]    reg_psum_15_23;
wire signed[15:0]    reg_weight_15_24;
wire signed[15:0]    reg_psum_15_24;
wire signed[15:0]    reg_weight_15_25;
wire signed[15:0]    reg_psum_15_25;
wire signed[15:0]    reg_weight_15_26;
wire signed[15:0]    reg_psum_15_26;
wire signed[15:0]    reg_weight_15_27;
wire signed[15:0]    reg_psum_15_27;
wire signed[15:0]    reg_weight_15_28;
wire signed[15:0]    reg_psum_15_28;
wire signed[15:0]    reg_weight_15_29;
wire signed[15:0]    reg_psum_15_29;
wire signed[15:0]    reg_weight_15_30;
wire signed[15:0]    reg_psum_15_30;
wire signed[15:0]    reg_weight_15_31;
wire signed[15:0]    reg_psum_15_31;
wire signed[15:0]    reg_weight_16_0;
wire signed[15:0]    reg_psum_16_0;
wire signed[15:0]    reg_weight_16_1;
wire signed[15:0]    reg_psum_16_1;
wire signed[15:0]    reg_weight_16_2;
wire signed[15:0]    reg_psum_16_2;
wire signed[15:0]    reg_weight_16_3;
wire signed[15:0]    reg_psum_16_3;
wire signed[15:0]    reg_weight_16_4;
wire signed[15:0]    reg_psum_16_4;
wire signed[15:0]    reg_weight_16_5;
wire signed[15:0]    reg_psum_16_5;
wire signed[15:0]    reg_weight_16_6;
wire signed[15:0]    reg_psum_16_6;
wire signed[15:0]    reg_weight_16_7;
wire signed[15:0]    reg_psum_16_7;
wire signed[15:0]    reg_weight_16_8;
wire signed[15:0]    reg_psum_16_8;
wire signed[15:0]    reg_weight_16_9;
wire signed[15:0]    reg_psum_16_9;
wire signed[15:0]    reg_weight_16_10;
wire signed[15:0]    reg_psum_16_10;
wire signed[15:0]    reg_weight_16_11;
wire signed[15:0]    reg_psum_16_11;
wire signed[15:0]    reg_weight_16_12;
wire signed[15:0]    reg_psum_16_12;
wire signed[15:0]    reg_weight_16_13;
wire signed[15:0]    reg_psum_16_13;
wire signed[15:0]    reg_weight_16_14;
wire signed[15:0]    reg_psum_16_14;
wire signed[15:0]    reg_weight_16_15;
wire signed[15:0]    reg_psum_16_15;
wire signed[15:0]    reg_weight_16_16;
wire signed[15:0]    reg_psum_16_16;
wire signed[15:0]    reg_weight_16_17;
wire signed[15:0]    reg_psum_16_17;
wire signed[15:0]    reg_weight_16_18;
wire signed[15:0]    reg_psum_16_18;
wire signed[15:0]    reg_weight_16_19;
wire signed[15:0]    reg_psum_16_19;
wire signed[15:0]    reg_weight_16_20;
wire signed[15:0]    reg_psum_16_20;
wire signed[15:0]    reg_weight_16_21;
wire signed[15:0]    reg_psum_16_21;
wire signed[15:0]    reg_weight_16_22;
wire signed[15:0]    reg_psum_16_22;
wire signed[15:0]    reg_weight_16_23;
wire signed[15:0]    reg_psum_16_23;
wire signed[15:0]    reg_weight_16_24;
wire signed[15:0]    reg_psum_16_24;
wire signed[15:0]    reg_weight_16_25;
wire signed[15:0]    reg_psum_16_25;
wire signed[15:0]    reg_weight_16_26;
wire signed[15:0]    reg_psum_16_26;
wire signed[15:0]    reg_weight_16_27;
wire signed[15:0]    reg_psum_16_27;
wire signed[15:0]    reg_weight_16_28;
wire signed[15:0]    reg_psum_16_28;
wire signed[15:0]    reg_weight_16_29;
wire signed[15:0]    reg_psum_16_29;
wire signed[15:0]    reg_weight_16_30;
wire signed[15:0]    reg_psum_16_30;
wire signed[15:0]    reg_weight_16_31;
wire signed[15:0]    reg_psum_16_31;
wire signed[15:0]    reg_weight_17_0;
wire signed[15:0]    reg_psum_17_0;
wire signed[15:0]    reg_weight_17_1;
wire signed[15:0]    reg_psum_17_1;
wire signed[15:0]    reg_weight_17_2;
wire signed[15:0]    reg_psum_17_2;
wire signed[15:0]    reg_weight_17_3;
wire signed[15:0]    reg_psum_17_3;
wire signed[15:0]    reg_weight_17_4;
wire signed[15:0]    reg_psum_17_4;
wire signed[15:0]    reg_weight_17_5;
wire signed[15:0]    reg_psum_17_5;
wire signed[15:0]    reg_weight_17_6;
wire signed[15:0]    reg_psum_17_6;
wire signed[15:0]    reg_weight_17_7;
wire signed[15:0]    reg_psum_17_7;
wire signed[15:0]    reg_weight_17_8;
wire signed[15:0]    reg_psum_17_8;
wire signed[15:0]    reg_weight_17_9;
wire signed[15:0]    reg_psum_17_9;
wire signed[15:0]    reg_weight_17_10;
wire signed[15:0]    reg_psum_17_10;
wire signed[15:0]    reg_weight_17_11;
wire signed[15:0]    reg_psum_17_11;
wire signed[15:0]    reg_weight_17_12;
wire signed[15:0]    reg_psum_17_12;
wire signed[15:0]    reg_weight_17_13;
wire signed[15:0]    reg_psum_17_13;
wire signed[15:0]    reg_weight_17_14;
wire signed[15:0]    reg_psum_17_14;
wire signed[15:0]    reg_weight_17_15;
wire signed[15:0]    reg_psum_17_15;
wire signed[15:0]    reg_weight_17_16;
wire signed[15:0]    reg_psum_17_16;
wire signed[15:0]    reg_weight_17_17;
wire signed[15:0]    reg_psum_17_17;
wire signed[15:0]    reg_weight_17_18;
wire signed[15:0]    reg_psum_17_18;
wire signed[15:0]    reg_weight_17_19;
wire signed[15:0]    reg_psum_17_19;
wire signed[15:0]    reg_weight_17_20;
wire signed[15:0]    reg_psum_17_20;
wire signed[15:0]    reg_weight_17_21;
wire signed[15:0]    reg_psum_17_21;
wire signed[15:0]    reg_weight_17_22;
wire signed[15:0]    reg_psum_17_22;
wire signed[15:0]    reg_weight_17_23;
wire signed[15:0]    reg_psum_17_23;
wire signed[15:0]    reg_weight_17_24;
wire signed[15:0]    reg_psum_17_24;
wire signed[15:0]    reg_weight_17_25;
wire signed[15:0]    reg_psum_17_25;
wire signed[15:0]    reg_weight_17_26;
wire signed[15:0]    reg_psum_17_26;
wire signed[15:0]    reg_weight_17_27;
wire signed[15:0]    reg_psum_17_27;
wire signed[15:0]    reg_weight_17_28;
wire signed[15:0]    reg_psum_17_28;
wire signed[15:0]    reg_weight_17_29;
wire signed[15:0]    reg_psum_17_29;
wire signed[15:0]    reg_weight_17_30;
wire signed[15:0]    reg_psum_17_30;
wire signed[15:0]    reg_weight_17_31;
wire signed[15:0]    reg_psum_17_31;
wire signed[15:0]    reg_weight_18_0;
wire signed[15:0]    reg_psum_18_0;
wire signed[15:0]    reg_weight_18_1;
wire signed[15:0]    reg_psum_18_1;
wire signed[15:0]    reg_weight_18_2;
wire signed[15:0]    reg_psum_18_2;
wire signed[15:0]    reg_weight_18_3;
wire signed[15:0]    reg_psum_18_3;
wire signed[15:0]    reg_weight_18_4;
wire signed[15:0]    reg_psum_18_4;
wire signed[15:0]    reg_weight_18_5;
wire signed[15:0]    reg_psum_18_5;
wire signed[15:0]    reg_weight_18_6;
wire signed[15:0]    reg_psum_18_6;
wire signed[15:0]    reg_weight_18_7;
wire signed[15:0]    reg_psum_18_7;
wire signed[15:0]    reg_weight_18_8;
wire signed[15:0]    reg_psum_18_8;
wire signed[15:0]    reg_weight_18_9;
wire signed[15:0]    reg_psum_18_9;
wire signed[15:0]    reg_weight_18_10;
wire signed[15:0]    reg_psum_18_10;
wire signed[15:0]    reg_weight_18_11;
wire signed[15:0]    reg_psum_18_11;
wire signed[15:0]    reg_weight_18_12;
wire signed[15:0]    reg_psum_18_12;
wire signed[15:0]    reg_weight_18_13;
wire signed[15:0]    reg_psum_18_13;
wire signed[15:0]    reg_weight_18_14;
wire signed[15:0]    reg_psum_18_14;
wire signed[15:0]    reg_weight_18_15;
wire signed[15:0]    reg_psum_18_15;
wire signed[15:0]    reg_weight_18_16;
wire signed[15:0]    reg_psum_18_16;
wire signed[15:0]    reg_weight_18_17;
wire signed[15:0]    reg_psum_18_17;
wire signed[15:0]    reg_weight_18_18;
wire signed[15:0]    reg_psum_18_18;
wire signed[15:0]    reg_weight_18_19;
wire signed[15:0]    reg_psum_18_19;
wire signed[15:0]    reg_weight_18_20;
wire signed[15:0]    reg_psum_18_20;
wire signed[15:0]    reg_weight_18_21;
wire signed[15:0]    reg_psum_18_21;
wire signed[15:0]    reg_weight_18_22;
wire signed[15:0]    reg_psum_18_22;
wire signed[15:0]    reg_weight_18_23;
wire signed[15:0]    reg_psum_18_23;
wire signed[15:0]    reg_weight_18_24;
wire signed[15:0]    reg_psum_18_24;
wire signed[15:0]    reg_weight_18_25;
wire signed[15:0]    reg_psum_18_25;
wire signed[15:0]    reg_weight_18_26;
wire signed[15:0]    reg_psum_18_26;
wire signed[15:0]    reg_weight_18_27;
wire signed[15:0]    reg_psum_18_27;
wire signed[15:0]    reg_weight_18_28;
wire signed[15:0]    reg_psum_18_28;
wire signed[15:0]    reg_weight_18_29;
wire signed[15:0]    reg_psum_18_29;
wire signed[15:0]    reg_weight_18_30;
wire signed[15:0]    reg_psum_18_30;
wire signed[15:0]    reg_weight_18_31;
wire signed[15:0]    reg_psum_18_31;
wire signed[15:0]    reg_weight_19_0;
wire signed[15:0]    reg_psum_19_0;
wire signed[15:0]    reg_weight_19_1;
wire signed[15:0]    reg_psum_19_1;
wire signed[15:0]    reg_weight_19_2;
wire signed[15:0]    reg_psum_19_2;
wire signed[15:0]    reg_weight_19_3;
wire signed[15:0]    reg_psum_19_3;
wire signed[15:0]    reg_weight_19_4;
wire signed[15:0]    reg_psum_19_4;
wire signed[15:0]    reg_weight_19_5;
wire signed[15:0]    reg_psum_19_5;
wire signed[15:0]    reg_weight_19_6;
wire signed[15:0]    reg_psum_19_6;
wire signed[15:0]    reg_weight_19_7;
wire signed[15:0]    reg_psum_19_7;
wire signed[15:0]    reg_weight_19_8;
wire signed[15:0]    reg_psum_19_8;
wire signed[15:0]    reg_weight_19_9;
wire signed[15:0]    reg_psum_19_9;
wire signed[15:0]    reg_weight_19_10;
wire signed[15:0]    reg_psum_19_10;
wire signed[15:0]    reg_weight_19_11;
wire signed[15:0]    reg_psum_19_11;
wire signed[15:0]    reg_weight_19_12;
wire signed[15:0]    reg_psum_19_12;
wire signed[15:0]    reg_weight_19_13;
wire signed[15:0]    reg_psum_19_13;
wire signed[15:0]    reg_weight_19_14;
wire signed[15:0]    reg_psum_19_14;
wire signed[15:0]    reg_weight_19_15;
wire signed[15:0]    reg_psum_19_15;
wire signed[15:0]    reg_weight_19_16;
wire signed[15:0]    reg_psum_19_16;
wire signed[15:0]    reg_weight_19_17;
wire signed[15:0]    reg_psum_19_17;
wire signed[15:0]    reg_weight_19_18;
wire signed[15:0]    reg_psum_19_18;
wire signed[15:0]    reg_weight_19_19;
wire signed[15:0]    reg_psum_19_19;
wire signed[15:0]    reg_weight_19_20;
wire signed[15:0]    reg_psum_19_20;
wire signed[15:0]    reg_weight_19_21;
wire signed[15:0]    reg_psum_19_21;
wire signed[15:0]    reg_weight_19_22;
wire signed[15:0]    reg_psum_19_22;
wire signed[15:0]    reg_weight_19_23;
wire signed[15:0]    reg_psum_19_23;
wire signed[15:0]    reg_weight_19_24;
wire signed[15:0]    reg_psum_19_24;
wire signed[15:0]    reg_weight_19_25;
wire signed[15:0]    reg_psum_19_25;
wire signed[15:0]    reg_weight_19_26;
wire signed[15:0]    reg_psum_19_26;
wire signed[15:0]    reg_weight_19_27;
wire signed[15:0]    reg_psum_19_27;
wire signed[15:0]    reg_weight_19_28;
wire signed[15:0]    reg_psum_19_28;
wire signed[15:0]    reg_weight_19_29;
wire signed[15:0]    reg_psum_19_29;
wire signed[15:0]    reg_weight_19_30;
wire signed[15:0]    reg_psum_19_30;
wire signed[15:0]    reg_weight_19_31;
wire signed[15:0]    reg_psum_19_31;
wire signed[15:0]    reg_weight_20_0;
wire signed[15:0]    reg_psum_20_0;
wire signed[15:0]    reg_weight_20_1;
wire signed[15:0]    reg_psum_20_1;
wire signed[15:0]    reg_weight_20_2;
wire signed[15:0]    reg_psum_20_2;
wire signed[15:0]    reg_weight_20_3;
wire signed[15:0]    reg_psum_20_3;
wire signed[15:0]    reg_weight_20_4;
wire signed[15:0]    reg_psum_20_4;
wire signed[15:0]    reg_weight_20_5;
wire signed[15:0]    reg_psum_20_5;
wire signed[15:0]    reg_weight_20_6;
wire signed[15:0]    reg_psum_20_6;
wire signed[15:0]    reg_weight_20_7;
wire signed[15:0]    reg_psum_20_7;
wire signed[15:0]    reg_weight_20_8;
wire signed[15:0]    reg_psum_20_8;
wire signed[15:0]    reg_weight_20_9;
wire signed[15:0]    reg_psum_20_9;
wire signed[15:0]    reg_weight_20_10;
wire signed[15:0]    reg_psum_20_10;
wire signed[15:0]    reg_weight_20_11;
wire signed[15:0]    reg_psum_20_11;
wire signed[15:0]    reg_weight_20_12;
wire signed[15:0]    reg_psum_20_12;
wire signed[15:0]    reg_weight_20_13;
wire signed[15:0]    reg_psum_20_13;
wire signed[15:0]    reg_weight_20_14;
wire signed[15:0]    reg_psum_20_14;
wire signed[15:0]    reg_weight_20_15;
wire signed[15:0]    reg_psum_20_15;
wire signed[15:0]    reg_weight_20_16;
wire signed[15:0]    reg_psum_20_16;
wire signed[15:0]    reg_weight_20_17;
wire signed[15:0]    reg_psum_20_17;
wire signed[15:0]    reg_weight_20_18;
wire signed[15:0]    reg_psum_20_18;
wire signed[15:0]    reg_weight_20_19;
wire signed[15:0]    reg_psum_20_19;
wire signed[15:0]    reg_weight_20_20;
wire signed[15:0]    reg_psum_20_20;
wire signed[15:0]    reg_weight_20_21;
wire signed[15:0]    reg_psum_20_21;
wire signed[15:0]    reg_weight_20_22;
wire signed[15:0]    reg_psum_20_22;
wire signed[15:0]    reg_weight_20_23;
wire signed[15:0]    reg_psum_20_23;
wire signed[15:0]    reg_weight_20_24;
wire signed[15:0]    reg_psum_20_24;
wire signed[15:0]    reg_weight_20_25;
wire signed[15:0]    reg_psum_20_25;
wire signed[15:0]    reg_weight_20_26;
wire signed[15:0]    reg_psum_20_26;
wire signed[15:0]    reg_weight_20_27;
wire signed[15:0]    reg_psum_20_27;
wire signed[15:0]    reg_weight_20_28;
wire signed[15:0]    reg_psum_20_28;
wire signed[15:0]    reg_weight_20_29;
wire signed[15:0]    reg_psum_20_29;
wire signed[15:0]    reg_weight_20_30;
wire signed[15:0]    reg_psum_20_30;
wire signed[15:0]    reg_weight_20_31;
wire signed[15:0]    reg_psum_20_31;
wire signed[15:0]    reg_weight_21_0;
wire signed[15:0]    reg_psum_21_0;
wire signed[15:0]    reg_weight_21_1;
wire signed[15:0]    reg_psum_21_1;
wire signed[15:0]    reg_weight_21_2;
wire signed[15:0]    reg_psum_21_2;
wire signed[15:0]    reg_weight_21_3;
wire signed[15:0]    reg_psum_21_3;
wire signed[15:0]    reg_weight_21_4;
wire signed[15:0]    reg_psum_21_4;
wire signed[15:0]    reg_weight_21_5;
wire signed[15:0]    reg_psum_21_5;
wire signed[15:0]    reg_weight_21_6;
wire signed[15:0]    reg_psum_21_6;
wire signed[15:0]    reg_weight_21_7;
wire signed[15:0]    reg_psum_21_7;
wire signed[15:0]    reg_weight_21_8;
wire signed[15:0]    reg_psum_21_8;
wire signed[15:0]    reg_weight_21_9;
wire signed[15:0]    reg_psum_21_9;
wire signed[15:0]    reg_weight_21_10;
wire signed[15:0]    reg_psum_21_10;
wire signed[15:0]    reg_weight_21_11;
wire signed[15:0]    reg_psum_21_11;
wire signed[15:0]    reg_weight_21_12;
wire signed[15:0]    reg_psum_21_12;
wire signed[15:0]    reg_weight_21_13;
wire signed[15:0]    reg_psum_21_13;
wire signed[15:0]    reg_weight_21_14;
wire signed[15:0]    reg_psum_21_14;
wire signed[15:0]    reg_weight_21_15;
wire signed[15:0]    reg_psum_21_15;
wire signed[15:0]    reg_weight_21_16;
wire signed[15:0]    reg_psum_21_16;
wire signed[15:0]    reg_weight_21_17;
wire signed[15:0]    reg_psum_21_17;
wire signed[15:0]    reg_weight_21_18;
wire signed[15:0]    reg_psum_21_18;
wire signed[15:0]    reg_weight_21_19;
wire signed[15:0]    reg_psum_21_19;
wire signed[15:0]    reg_weight_21_20;
wire signed[15:0]    reg_psum_21_20;
wire signed[15:0]    reg_weight_21_21;
wire signed[15:0]    reg_psum_21_21;
wire signed[15:0]    reg_weight_21_22;
wire signed[15:0]    reg_psum_21_22;
wire signed[15:0]    reg_weight_21_23;
wire signed[15:0]    reg_psum_21_23;
wire signed[15:0]    reg_weight_21_24;
wire signed[15:0]    reg_psum_21_24;
wire signed[15:0]    reg_weight_21_25;
wire signed[15:0]    reg_psum_21_25;
wire signed[15:0]    reg_weight_21_26;
wire signed[15:0]    reg_psum_21_26;
wire signed[15:0]    reg_weight_21_27;
wire signed[15:0]    reg_psum_21_27;
wire signed[15:0]    reg_weight_21_28;
wire signed[15:0]    reg_psum_21_28;
wire signed[15:0]    reg_weight_21_29;
wire signed[15:0]    reg_psum_21_29;
wire signed[15:0]    reg_weight_21_30;
wire signed[15:0]    reg_psum_21_30;
wire signed[15:0]    reg_weight_21_31;
wire signed[15:0]    reg_psum_21_31;
wire signed[15:0]    reg_weight_22_0;
wire signed[15:0]    reg_psum_22_0;
wire signed[15:0]    reg_weight_22_1;
wire signed[15:0]    reg_psum_22_1;
wire signed[15:0]    reg_weight_22_2;
wire signed[15:0]    reg_psum_22_2;
wire signed[15:0]    reg_weight_22_3;
wire signed[15:0]    reg_psum_22_3;
wire signed[15:0]    reg_weight_22_4;
wire signed[15:0]    reg_psum_22_4;
wire signed[15:0]    reg_weight_22_5;
wire signed[15:0]    reg_psum_22_5;
wire signed[15:0]    reg_weight_22_6;
wire signed[15:0]    reg_psum_22_6;
wire signed[15:0]    reg_weight_22_7;
wire signed[15:0]    reg_psum_22_7;
wire signed[15:0]    reg_weight_22_8;
wire signed[15:0]    reg_psum_22_8;
wire signed[15:0]    reg_weight_22_9;
wire signed[15:0]    reg_psum_22_9;
wire signed[15:0]    reg_weight_22_10;
wire signed[15:0]    reg_psum_22_10;
wire signed[15:0]    reg_weight_22_11;
wire signed[15:0]    reg_psum_22_11;
wire signed[15:0]    reg_weight_22_12;
wire signed[15:0]    reg_psum_22_12;
wire signed[15:0]    reg_weight_22_13;
wire signed[15:0]    reg_psum_22_13;
wire signed[15:0]    reg_weight_22_14;
wire signed[15:0]    reg_psum_22_14;
wire signed[15:0]    reg_weight_22_15;
wire signed[15:0]    reg_psum_22_15;
wire signed[15:0]    reg_weight_22_16;
wire signed[15:0]    reg_psum_22_16;
wire signed[15:0]    reg_weight_22_17;
wire signed[15:0]    reg_psum_22_17;
wire signed[15:0]    reg_weight_22_18;
wire signed[15:0]    reg_psum_22_18;
wire signed[15:0]    reg_weight_22_19;
wire signed[15:0]    reg_psum_22_19;
wire signed[15:0]    reg_weight_22_20;
wire signed[15:0]    reg_psum_22_20;
wire signed[15:0]    reg_weight_22_21;
wire signed[15:0]    reg_psum_22_21;
wire signed[15:0]    reg_weight_22_22;
wire signed[15:0]    reg_psum_22_22;
wire signed[15:0]    reg_weight_22_23;
wire signed[15:0]    reg_psum_22_23;
wire signed[15:0]    reg_weight_22_24;
wire signed[15:0]    reg_psum_22_24;
wire signed[15:0]    reg_weight_22_25;
wire signed[15:0]    reg_psum_22_25;
wire signed[15:0]    reg_weight_22_26;
wire signed[15:0]    reg_psum_22_26;
wire signed[15:0]    reg_weight_22_27;
wire signed[15:0]    reg_psum_22_27;
wire signed[15:0]    reg_weight_22_28;
wire signed[15:0]    reg_psum_22_28;
wire signed[15:0]    reg_weight_22_29;
wire signed[15:0]    reg_psum_22_29;
wire signed[15:0]    reg_weight_22_30;
wire signed[15:0]    reg_psum_22_30;
wire signed[15:0]    reg_weight_22_31;
wire signed[15:0]    reg_psum_22_31;
wire signed[15:0]    reg_weight_23_0;
wire signed[15:0]    reg_psum_23_0;
wire signed[15:0]    reg_weight_23_1;
wire signed[15:0]    reg_psum_23_1;
wire signed[15:0]    reg_weight_23_2;
wire signed[15:0]    reg_psum_23_2;
wire signed[15:0]    reg_weight_23_3;
wire signed[15:0]    reg_psum_23_3;
wire signed[15:0]    reg_weight_23_4;
wire signed[15:0]    reg_psum_23_4;
wire signed[15:0]    reg_weight_23_5;
wire signed[15:0]    reg_psum_23_5;
wire signed[15:0]    reg_weight_23_6;
wire signed[15:0]    reg_psum_23_6;
wire signed[15:0]    reg_weight_23_7;
wire signed[15:0]    reg_psum_23_7;
wire signed[15:0]    reg_weight_23_8;
wire signed[15:0]    reg_psum_23_8;
wire signed[15:0]    reg_weight_23_9;
wire signed[15:0]    reg_psum_23_9;
wire signed[15:0]    reg_weight_23_10;
wire signed[15:0]    reg_psum_23_10;
wire signed[15:0]    reg_weight_23_11;
wire signed[15:0]    reg_psum_23_11;
wire signed[15:0]    reg_weight_23_12;
wire signed[15:0]    reg_psum_23_12;
wire signed[15:0]    reg_weight_23_13;
wire signed[15:0]    reg_psum_23_13;
wire signed[15:0]    reg_weight_23_14;
wire signed[15:0]    reg_psum_23_14;
wire signed[15:0]    reg_weight_23_15;
wire signed[15:0]    reg_psum_23_15;
wire signed[15:0]    reg_weight_23_16;
wire signed[15:0]    reg_psum_23_16;
wire signed[15:0]    reg_weight_23_17;
wire signed[15:0]    reg_psum_23_17;
wire signed[15:0]    reg_weight_23_18;
wire signed[15:0]    reg_psum_23_18;
wire signed[15:0]    reg_weight_23_19;
wire signed[15:0]    reg_psum_23_19;
wire signed[15:0]    reg_weight_23_20;
wire signed[15:0]    reg_psum_23_20;
wire signed[15:0]    reg_weight_23_21;
wire signed[15:0]    reg_psum_23_21;
wire signed[15:0]    reg_weight_23_22;
wire signed[15:0]    reg_psum_23_22;
wire signed[15:0]    reg_weight_23_23;
wire signed[15:0]    reg_psum_23_23;
wire signed[15:0]    reg_weight_23_24;
wire signed[15:0]    reg_psum_23_24;
wire signed[15:0]    reg_weight_23_25;
wire signed[15:0]    reg_psum_23_25;
wire signed[15:0]    reg_weight_23_26;
wire signed[15:0]    reg_psum_23_26;
wire signed[15:0]    reg_weight_23_27;
wire signed[15:0]    reg_psum_23_27;
wire signed[15:0]    reg_weight_23_28;
wire signed[15:0]    reg_psum_23_28;
wire signed[15:0]    reg_weight_23_29;
wire signed[15:0]    reg_psum_23_29;
wire signed[15:0]    reg_weight_23_30;
wire signed[15:0]    reg_psum_23_30;
wire signed[15:0]    reg_weight_23_31;
wire signed[15:0]    reg_psum_23_31;
wire signed[15:0]    reg_weight_24_0;
wire signed[15:0]    reg_psum_24_0;
wire signed[15:0]    reg_weight_24_1;
wire signed[15:0]    reg_psum_24_1;
wire signed[15:0]    reg_weight_24_2;
wire signed[15:0]    reg_psum_24_2;
wire signed[15:0]    reg_weight_24_3;
wire signed[15:0]    reg_psum_24_3;
wire signed[15:0]    reg_weight_24_4;
wire signed[15:0]    reg_psum_24_4;
wire signed[15:0]    reg_weight_24_5;
wire signed[15:0]    reg_psum_24_5;
wire signed[15:0]    reg_weight_24_6;
wire signed[15:0]    reg_psum_24_6;
wire signed[15:0]    reg_weight_24_7;
wire signed[15:0]    reg_psum_24_7;
wire signed[15:0]    reg_weight_24_8;
wire signed[15:0]    reg_psum_24_8;
wire signed[15:0]    reg_weight_24_9;
wire signed[15:0]    reg_psum_24_9;
wire signed[15:0]    reg_weight_24_10;
wire signed[15:0]    reg_psum_24_10;
wire signed[15:0]    reg_weight_24_11;
wire signed[15:0]    reg_psum_24_11;
wire signed[15:0]    reg_weight_24_12;
wire signed[15:0]    reg_psum_24_12;
wire signed[15:0]    reg_weight_24_13;
wire signed[15:0]    reg_psum_24_13;
wire signed[15:0]    reg_weight_24_14;
wire signed[15:0]    reg_psum_24_14;
wire signed[15:0]    reg_weight_24_15;
wire signed[15:0]    reg_psum_24_15;
wire signed[15:0]    reg_weight_24_16;
wire signed[15:0]    reg_psum_24_16;
wire signed[15:0]    reg_weight_24_17;
wire signed[15:0]    reg_psum_24_17;
wire signed[15:0]    reg_weight_24_18;
wire signed[15:0]    reg_psum_24_18;
wire signed[15:0]    reg_weight_24_19;
wire signed[15:0]    reg_psum_24_19;
wire signed[15:0]    reg_weight_24_20;
wire signed[15:0]    reg_psum_24_20;
wire signed[15:0]    reg_weight_24_21;
wire signed[15:0]    reg_psum_24_21;
wire signed[15:0]    reg_weight_24_22;
wire signed[15:0]    reg_psum_24_22;
wire signed[15:0]    reg_weight_24_23;
wire signed[15:0]    reg_psum_24_23;
wire signed[15:0]    reg_weight_24_24;
wire signed[15:0]    reg_psum_24_24;
wire signed[15:0]    reg_weight_24_25;
wire signed[15:0]    reg_psum_24_25;
wire signed[15:0]    reg_weight_24_26;
wire signed[15:0]    reg_psum_24_26;
wire signed[15:0]    reg_weight_24_27;
wire signed[15:0]    reg_psum_24_27;
wire signed[15:0]    reg_weight_24_28;
wire signed[15:0]    reg_psum_24_28;
wire signed[15:0]    reg_weight_24_29;
wire signed[15:0]    reg_psum_24_29;
wire signed[15:0]    reg_weight_24_30;
wire signed[15:0]    reg_psum_24_30;
wire signed[15:0]    reg_weight_24_31;
wire signed[15:0]    reg_psum_24_31;
wire signed[15:0]    reg_weight_25_0;
wire signed[15:0]    reg_psum_25_0;
wire signed[15:0]    reg_weight_25_1;
wire signed[15:0]    reg_psum_25_1;
wire signed[15:0]    reg_weight_25_2;
wire signed[15:0]    reg_psum_25_2;
wire signed[15:0]    reg_weight_25_3;
wire signed[15:0]    reg_psum_25_3;
wire signed[15:0]    reg_weight_25_4;
wire signed[15:0]    reg_psum_25_4;
wire signed[15:0]    reg_weight_25_5;
wire signed[15:0]    reg_psum_25_5;
wire signed[15:0]    reg_weight_25_6;
wire signed[15:0]    reg_psum_25_6;
wire signed[15:0]    reg_weight_25_7;
wire signed[15:0]    reg_psum_25_7;
wire signed[15:0]    reg_weight_25_8;
wire signed[15:0]    reg_psum_25_8;
wire signed[15:0]    reg_weight_25_9;
wire signed[15:0]    reg_psum_25_9;
wire signed[15:0]    reg_weight_25_10;
wire signed[15:0]    reg_psum_25_10;
wire signed[15:0]    reg_weight_25_11;
wire signed[15:0]    reg_psum_25_11;
wire signed[15:0]    reg_weight_25_12;
wire signed[15:0]    reg_psum_25_12;
wire signed[15:0]    reg_weight_25_13;
wire signed[15:0]    reg_psum_25_13;
wire signed[15:0]    reg_weight_25_14;
wire signed[15:0]    reg_psum_25_14;
wire signed[15:0]    reg_weight_25_15;
wire signed[15:0]    reg_psum_25_15;
wire signed[15:0]    reg_weight_25_16;
wire signed[15:0]    reg_psum_25_16;
wire signed[15:0]    reg_weight_25_17;
wire signed[15:0]    reg_psum_25_17;
wire signed[15:0]    reg_weight_25_18;
wire signed[15:0]    reg_psum_25_18;
wire signed[15:0]    reg_weight_25_19;
wire signed[15:0]    reg_psum_25_19;
wire signed[15:0]    reg_weight_25_20;
wire signed[15:0]    reg_psum_25_20;
wire signed[15:0]    reg_weight_25_21;
wire signed[15:0]    reg_psum_25_21;
wire signed[15:0]    reg_weight_25_22;
wire signed[15:0]    reg_psum_25_22;
wire signed[15:0]    reg_weight_25_23;
wire signed[15:0]    reg_psum_25_23;
wire signed[15:0]    reg_weight_25_24;
wire signed[15:0]    reg_psum_25_24;
wire signed[15:0]    reg_weight_25_25;
wire signed[15:0]    reg_psum_25_25;
wire signed[15:0]    reg_weight_25_26;
wire signed[15:0]    reg_psum_25_26;
wire signed[15:0]    reg_weight_25_27;
wire signed[15:0]    reg_psum_25_27;
wire signed[15:0]    reg_weight_25_28;
wire signed[15:0]    reg_psum_25_28;
wire signed[15:0]    reg_weight_25_29;
wire signed[15:0]    reg_psum_25_29;
wire signed[15:0]    reg_weight_25_30;
wire signed[15:0]    reg_psum_25_30;
wire signed[15:0]    reg_weight_25_31;
wire signed[15:0]    reg_psum_25_31;
wire signed[15:0]    reg_weight_26_0;
wire signed[15:0]    reg_psum_26_0;
wire signed[15:0]    reg_weight_26_1;
wire signed[15:0]    reg_psum_26_1;
wire signed[15:0]    reg_weight_26_2;
wire signed[15:0]    reg_psum_26_2;
wire signed[15:0]    reg_weight_26_3;
wire signed[15:0]    reg_psum_26_3;
wire signed[15:0]    reg_weight_26_4;
wire signed[15:0]    reg_psum_26_4;
wire signed[15:0]    reg_weight_26_5;
wire signed[15:0]    reg_psum_26_5;
wire signed[15:0]    reg_weight_26_6;
wire signed[15:0]    reg_psum_26_6;
wire signed[15:0]    reg_weight_26_7;
wire signed[15:0]    reg_psum_26_7;
wire signed[15:0]    reg_weight_26_8;
wire signed[15:0]    reg_psum_26_8;
wire signed[15:0]    reg_weight_26_9;
wire signed[15:0]    reg_psum_26_9;
wire signed[15:0]    reg_weight_26_10;
wire signed[15:0]    reg_psum_26_10;
wire signed[15:0]    reg_weight_26_11;
wire signed[15:0]    reg_psum_26_11;
wire signed[15:0]    reg_weight_26_12;
wire signed[15:0]    reg_psum_26_12;
wire signed[15:0]    reg_weight_26_13;
wire signed[15:0]    reg_psum_26_13;
wire signed[15:0]    reg_weight_26_14;
wire signed[15:0]    reg_psum_26_14;
wire signed[15:0]    reg_weight_26_15;
wire signed[15:0]    reg_psum_26_15;
wire signed[15:0]    reg_weight_26_16;
wire signed[15:0]    reg_psum_26_16;
wire signed[15:0]    reg_weight_26_17;
wire signed[15:0]    reg_psum_26_17;
wire signed[15:0]    reg_weight_26_18;
wire signed[15:0]    reg_psum_26_18;
wire signed[15:0]    reg_weight_26_19;
wire signed[15:0]    reg_psum_26_19;
wire signed[15:0]    reg_weight_26_20;
wire signed[15:0]    reg_psum_26_20;
wire signed[15:0]    reg_weight_26_21;
wire signed[15:0]    reg_psum_26_21;
wire signed[15:0]    reg_weight_26_22;
wire signed[15:0]    reg_psum_26_22;
wire signed[15:0]    reg_weight_26_23;
wire signed[15:0]    reg_psum_26_23;
wire signed[15:0]    reg_weight_26_24;
wire signed[15:0]    reg_psum_26_24;
wire signed[15:0]    reg_weight_26_25;
wire signed[15:0]    reg_psum_26_25;
wire signed[15:0]    reg_weight_26_26;
wire signed[15:0]    reg_psum_26_26;
wire signed[15:0]    reg_weight_26_27;
wire signed[15:0]    reg_psum_26_27;
wire signed[15:0]    reg_weight_26_28;
wire signed[15:0]    reg_psum_26_28;
wire signed[15:0]    reg_weight_26_29;
wire signed[15:0]    reg_psum_26_29;
wire signed[15:0]    reg_weight_26_30;
wire signed[15:0]    reg_psum_26_30;
wire signed[15:0]    reg_weight_26_31;
wire signed[15:0]    reg_psum_26_31;
wire signed[15:0]    reg_weight_27_0;
wire signed[15:0]    reg_psum_27_0;
wire signed[15:0]    reg_weight_27_1;
wire signed[15:0]    reg_psum_27_1;
wire signed[15:0]    reg_weight_27_2;
wire signed[15:0]    reg_psum_27_2;
wire signed[15:0]    reg_weight_27_3;
wire signed[15:0]    reg_psum_27_3;
wire signed[15:0]    reg_weight_27_4;
wire signed[15:0]    reg_psum_27_4;
wire signed[15:0]    reg_weight_27_5;
wire signed[15:0]    reg_psum_27_5;
wire signed[15:0]    reg_weight_27_6;
wire signed[15:0]    reg_psum_27_6;
wire signed[15:0]    reg_weight_27_7;
wire signed[15:0]    reg_psum_27_7;
wire signed[15:0]    reg_weight_27_8;
wire signed[15:0]    reg_psum_27_8;
wire signed[15:0]    reg_weight_27_9;
wire signed[15:0]    reg_psum_27_9;
wire signed[15:0]    reg_weight_27_10;
wire signed[15:0]    reg_psum_27_10;
wire signed[15:0]    reg_weight_27_11;
wire signed[15:0]    reg_psum_27_11;
wire signed[15:0]    reg_weight_27_12;
wire signed[15:0]    reg_psum_27_12;
wire signed[15:0]    reg_weight_27_13;
wire signed[15:0]    reg_psum_27_13;
wire signed[15:0]    reg_weight_27_14;
wire signed[15:0]    reg_psum_27_14;
wire signed[15:0]    reg_weight_27_15;
wire signed[15:0]    reg_psum_27_15;
wire signed[15:0]    reg_weight_27_16;
wire signed[15:0]    reg_psum_27_16;
wire signed[15:0]    reg_weight_27_17;
wire signed[15:0]    reg_psum_27_17;
wire signed[15:0]    reg_weight_27_18;
wire signed[15:0]    reg_psum_27_18;
wire signed[15:0]    reg_weight_27_19;
wire signed[15:0]    reg_psum_27_19;
wire signed[15:0]    reg_weight_27_20;
wire signed[15:0]    reg_psum_27_20;
wire signed[15:0]    reg_weight_27_21;
wire signed[15:0]    reg_psum_27_21;
wire signed[15:0]    reg_weight_27_22;
wire signed[15:0]    reg_psum_27_22;
wire signed[15:0]    reg_weight_27_23;
wire signed[15:0]    reg_psum_27_23;
wire signed[15:0]    reg_weight_27_24;
wire signed[15:0]    reg_psum_27_24;
wire signed[15:0]    reg_weight_27_25;
wire signed[15:0]    reg_psum_27_25;
wire signed[15:0]    reg_weight_27_26;
wire signed[15:0]    reg_psum_27_26;
wire signed[15:0]    reg_weight_27_27;
wire signed[15:0]    reg_psum_27_27;
wire signed[15:0]    reg_weight_27_28;
wire signed[15:0]    reg_psum_27_28;
wire signed[15:0]    reg_weight_27_29;
wire signed[15:0]    reg_psum_27_29;
wire signed[15:0]    reg_weight_27_30;
wire signed[15:0]    reg_psum_27_30;
wire signed[15:0]    reg_weight_27_31;
wire signed[15:0]    reg_psum_27_31;
wire signed[15:0]    reg_weight_28_0;
wire signed[15:0]    reg_psum_28_0;
wire signed[15:0]    reg_weight_28_1;
wire signed[15:0]    reg_psum_28_1;
wire signed[15:0]    reg_weight_28_2;
wire signed[15:0]    reg_psum_28_2;
wire signed[15:0]    reg_weight_28_3;
wire signed[15:0]    reg_psum_28_3;
wire signed[15:0]    reg_weight_28_4;
wire signed[15:0]    reg_psum_28_4;
wire signed[15:0]    reg_weight_28_5;
wire signed[15:0]    reg_psum_28_5;
wire signed[15:0]    reg_weight_28_6;
wire signed[15:0]    reg_psum_28_6;
wire signed[15:0]    reg_weight_28_7;
wire signed[15:0]    reg_psum_28_7;
wire signed[15:0]    reg_weight_28_8;
wire signed[15:0]    reg_psum_28_8;
wire signed[15:0]    reg_weight_28_9;
wire signed[15:0]    reg_psum_28_9;
wire signed[15:0]    reg_weight_28_10;
wire signed[15:0]    reg_psum_28_10;
wire signed[15:0]    reg_weight_28_11;
wire signed[15:0]    reg_psum_28_11;
wire signed[15:0]    reg_weight_28_12;
wire signed[15:0]    reg_psum_28_12;
wire signed[15:0]    reg_weight_28_13;
wire signed[15:0]    reg_psum_28_13;
wire signed[15:0]    reg_weight_28_14;
wire signed[15:0]    reg_psum_28_14;
wire signed[15:0]    reg_weight_28_15;
wire signed[15:0]    reg_psum_28_15;
wire signed[15:0]    reg_weight_28_16;
wire signed[15:0]    reg_psum_28_16;
wire signed[15:0]    reg_weight_28_17;
wire signed[15:0]    reg_psum_28_17;
wire signed[15:0]    reg_weight_28_18;
wire signed[15:0]    reg_psum_28_18;
wire signed[15:0]    reg_weight_28_19;
wire signed[15:0]    reg_psum_28_19;
wire signed[15:0]    reg_weight_28_20;
wire signed[15:0]    reg_psum_28_20;
wire signed[15:0]    reg_weight_28_21;
wire signed[15:0]    reg_psum_28_21;
wire signed[15:0]    reg_weight_28_22;
wire signed[15:0]    reg_psum_28_22;
wire signed[15:0]    reg_weight_28_23;
wire signed[15:0]    reg_psum_28_23;
wire signed[15:0]    reg_weight_28_24;
wire signed[15:0]    reg_psum_28_24;
wire signed[15:0]    reg_weight_28_25;
wire signed[15:0]    reg_psum_28_25;
wire signed[15:0]    reg_weight_28_26;
wire signed[15:0]    reg_psum_28_26;
wire signed[15:0]    reg_weight_28_27;
wire signed[15:0]    reg_psum_28_27;
wire signed[15:0]    reg_weight_28_28;
wire signed[15:0]    reg_psum_28_28;
wire signed[15:0]    reg_weight_28_29;
wire signed[15:0]    reg_psum_28_29;
wire signed[15:0]    reg_weight_28_30;
wire signed[15:0]    reg_psum_28_30;
wire signed[15:0]    reg_weight_28_31;
wire signed[15:0]    reg_psum_28_31;
wire signed[15:0]    reg_weight_29_0;
wire signed[15:0]    reg_psum_29_0;
wire signed[15:0]    reg_weight_29_1;
wire signed[15:0]    reg_psum_29_1;
wire signed[15:0]    reg_weight_29_2;
wire signed[15:0]    reg_psum_29_2;
wire signed[15:0]    reg_weight_29_3;
wire signed[15:0]    reg_psum_29_3;
wire signed[15:0]    reg_weight_29_4;
wire signed[15:0]    reg_psum_29_4;
wire signed[15:0]    reg_weight_29_5;
wire signed[15:0]    reg_psum_29_5;
wire signed[15:0]    reg_weight_29_6;
wire signed[15:0]    reg_psum_29_6;
wire signed[15:0]    reg_weight_29_7;
wire signed[15:0]    reg_psum_29_7;
wire signed[15:0]    reg_weight_29_8;
wire signed[15:0]    reg_psum_29_8;
wire signed[15:0]    reg_weight_29_9;
wire signed[15:0]    reg_psum_29_9;
wire signed[15:0]    reg_weight_29_10;
wire signed[15:0]    reg_psum_29_10;
wire signed[15:0]    reg_weight_29_11;
wire signed[15:0]    reg_psum_29_11;
wire signed[15:0]    reg_weight_29_12;
wire signed[15:0]    reg_psum_29_12;
wire signed[15:0]    reg_weight_29_13;
wire signed[15:0]    reg_psum_29_13;
wire signed[15:0]    reg_weight_29_14;
wire signed[15:0]    reg_psum_29_14;
wire signed[15:0]    reg_weight_29_15;
wire signed[15:0]    reg_psum_29_15;
wire signed[15:0]    reg_weight_29_16;
wire signed[15:0]    reg_psum_29_16;
wire signed[15:0]    reg_weight_29_17;
wire signed[15:0]    reg_psum_29_17;
wire signed[15:0]    reg_weight_29_18;
wire signed[15:0]    reg_psum_29_18;
wire signed[15:0]    reg_weight_29_19;
wire signed[15:0]    reg_psum_29_19;
wire signed[15:0]    reg_weight_29_20;
wire signed[15:0]    reg_psum_29_20;
wire signed[15:0]    reg_weight_29_21;
wire signed[15:0]    reg_psum_29_21;
wire signed[15:0]    reg_weight_29_22;
wire signed[15:0]    reg_psum_29_22;
wire signed[15:0]    reg_weight_29_23;
wire signed[15:0]    reg_psum_29_23;
wire signed[15:0]    reg_weight_29_24;
wire signed[15:0]    reg_psum_29_24;
wire signed[15:0]    reg_weight_29_25;
wire signed[15:0]    reg_psum_29_25;
wire signed[15:0]    reg_weight_29_26;
wire signed[15:0]    reg_psum_29_26;
wire signed[15:0]    reg_weight_29_27;
wire signed[15:0]    reg_psum_29_27;
wire signed[15:0]    reg_weight_29_28;
wire signed[15:0]    reg_psum_29_28;
wire signed[15:0]    reg_weight_29_29;
wire signed[15:0]    reg_psum_29_29;
wire signed[15:0]    reg_weight_29_30;
wire signed[15:0]    reg_psum_29_30;
wire signed[15:0]    reg_weight_29_31;
wire signed[15:0]    reg_psum_29_31;
wire signed[15:0]    reg_weight_30_0;
wire signed[15:0]    reg_psum_30_0;
wire signed[15:0]    reg_weight_30_1;
wire signed[15:0]    reg_psum_30_1;
wire signed[15:0]    reg_weight_30_2;
wire signed[15:0]    reg_psum_30_2;
wire signed[15:0]    reg_weight_30_3;
wire signed[15:0]    reg_psum_30_3;
wire signed[15:0]    reg_weight_30_4;
wire signed[15:0]    reg_psum_30_4;
wire signed[15:0]    reg_weight_30_5;
wire signed[15:0]    reg_psum_30_5;
wire signed[15:0]    reg_weight_30_6;
wire signed[15:0]    reg_psum_30_6;
wire signed[15:0]    reg_weight_30_7;
wire signed[15:0]    reg_psum_30_7;
wire signed[15:0]    reg_weight_30_8;
wire signed[15:0]    reg_psum_30_8;
wire signed[15:0]    reg_weight_30_9;
wire signed[15:0]    reg_psum_30_9;
wire signed[15:0]    reg_weight_30_10;
wire signed[15:0]    reg_psum_30_10;
wire signed[15:0]    reg_weight_30_11;
wire signed[15:0]    reg_psum_30_11;
wire signed[15:0]    reg_weight_30_12;
wire signed[15:0]    reg_psum_30_12;
wire signed[15:0]    reg_weight_30_13;
wire signed[15:0]    reg_psum_30_13;
wire signed[15:0]    reg_weight_30_14;
wire signed[15:0]    reg_psum_30_14;
wire signed[15:0]    reg_weight_30_15;
wire signed[15:0]    reg_psum_30_15;
wire signed[15:0]    reg_weight_30_16;
wire signed[15:0]    reg_psum_30_16;
wire signed[15:0]    reg_weight_30_17;
wire signed[15:0]    reg_psum_30_17;
wire signed[15:0]    reg_weight_30_18;
wire signed[15:0]    reg_psum_30_18;
wire signed[15:0]    reg_weight_30_19;
wire signed[15:0]    reg_psum_30_19;
wire signed[15:0]    reg_weight_30_20;
wire signed[15:0]    reg_psum_30_20;
wire signed[15:0]    reg_weight_30_21;
wire signed[15:0]    reg_psum_30_21;
wire signed[15:0]    reg_weight_30_22;
wire signed[15:0]    reg_psum_30_22;
wire signed[15:0]    reg_weight_30_23;
wire signed[15:0]    reg_psum_30_23;
wire signed[15:0]    reg_weight_30_24;
wire signed[15:0]    reg_psum_30_24;
wire signed[15:0]    reg_weight_30_25;
wire signed[15:0]    reg_psum_30_25;
wire signed[15:0]    reg_weight_30_26;
wire signed[15:0]    reg_psum_30_26;
wire signed[15:0]    reg_weight_30_27;
wire signed[15:0]    reg_psum_30_27;
wire signed[15:0]    reg_weight_30_28;
wire signed[15:0]    reg_psum_30_28;
wire signed[15:0]    reg_weight_30_29;
wire signed[15:0]    reg_psum_30_29;
wire signed[15:0]    reg_weight_30_30;
wire signed[15:0]    reg_psum_30_30;
wire signed[15:0]    reg_weight_30_31;
wire signed[15:0]    reg_psum_30_31;
wire signed[15:0]    reg_weight_31_0;
wire signed[15:0]    reg_psum_31_0;
wire signed[15:0]    reg_weight_31_1;
wire signed[15:0]    reg_psum_31_1;
wire signed[15:0]    reg_weight_31_2;
wire signed[15:0]    reg_psum_31_2;
wire signed[15:0]    reg_weight_31_3;
wire signed[15:0]    reg_psum_31_3;
wire signed[15:0]    reg_weight_31_4;
wire signed[15:0]    reg_psum_31_4;
wire signed[15:0]    reg_weight_31_5;
wire signed[15:0]    reg_psum_31_5;
wire signed[15:0]    reg_weight_31_6;
wire signed[15:0]    reg_psum_31_6;
wire signed[15:0]    reg_weight_31_7;
wire signed[15:0]    reg_psum_31_7;
wire signed[15:0]    reg_weight_31_8;
wire signed[15:0]    reg_psum_31_8;
wire signed[15:0]    reg_weight_31_9;
wire signed[15:0]    reg_psum_31_9;
wire signed[15:0]    reg_weight_31_10;
wire signed[15:0]    reg_psum_31_10;
wire signed[15:0]    reg_weight_31_11;
wire signed[15:0]    reg_psum_31_11;
wire signed[15:0]    reg_weight_31_12;
wire signed[15:0]    reg_psum_31_12;
wire signed[15:0]    reg_weight_31_13;
wire signed[15:0]    reg_psum_31_13;
wire signed[15:0]    reg_weight_31_14;
wire signed[15:0]    reg_psum_31_14;
wire signed[15:0]    reg_weight_31_15;
wire signed[15:0]    reg_psum_31_15;
wire signed[15:0]    reg_weight_31_16;
wire signed[15:0]    reg_psum_31_16;
wire signed[15:0]    reg_weight_31_17;
wire signed[15:0]    reg_psum_31_17;
wire signed[15:0]    reg_weight_31_18;
wire signed[15:0]    reg_psum_31_18;
wire signed[15:0]    reg_weight_31_19;
wire signed[15:0]    reg_psum_31_19;
wire signed[15:0]    reg_weight_31_20;
wire signed[15:0]    reg_psum_31_20;
wire signed[15:0]    reg_weight_31_21;
wire signed[15:0]    reg_psum_31_21;
wire signed[15:0]    reg_weight_31_22;
wire signed[15:0]    reg_psum_31_22;
wire signed[15:0]    reg_weight_31_23;
wire signed[15:0]    reg_psum_31_23;
wire signed[15:0]    reg_weight_31_24;
wire signed[15:0]    reg_psum_31_24;
wire signed[15:0]    reg_weight_31_25;
wire signed[15:0]    reg_psum_31_25;
wire signed[15:0]    reg_weight_31_26;
wire signed[15:0]    reg_psum_31_26;
wire signed[15:0]    reg_weight_31_27;
wire signed[15:0]    reg_psum_31_27;
wire signed[15:0]    reg_weight_31_28;
wire signed[15:0]    reg_psum_31_28;
wire signed[15:0]    reg_weight_31_29;
wire signed[15:0]    reg_psum_31_29;
wire signed[15:0]    reg_weight_31_30;
wire signed[15:0]    reg_psum_31_30;
wire signed[15:0]    reg_weight_31_31;
wire signed[15:0]    reg_psum_31_31;
assign out_psum_0 =  reg_psum_31_0;
assign out_psum_1 =  reg_psum_31_1;
assign out_psum_2 =  reg_psum_31_2;
assign out_psum_3 =  reg_psum_31_3;
assign out_psum_4 =  reg_psum_31_4;
assign out_psum_5 =  reg_psum_31_5;
assign out_psum_6 =  reg_psum_31_6;
assign out_psum_7 =  reg_psum_31_7;
assign out_psum_8 =  reg_psum_31_8;
assign out_psum_9 =  reg_psum_31_9;
assign out_psum_10 =  reg_psum_31_10;
assign out_psum_11 =  reg_psum_31_11;
assign out_psum_12 =  reg_psum_31_12;
assign out_psum_13 =  reg_psum_31_13;
assign out_psum_14 =  reg_psum_31_14;
assign out_psum_15 =  reg_psum_31_15;
assign out_psum_16 =  reg_psum_31_16;
assign out_psum_17 =  reg_psum_31_17;
assign out_psum_18 =  reg_psum_31_18;
assign out_psum_19 =  reg_psum_31_19;
assign out_psum_20 =  reg_psum_31_20;
assign out_psum_21 =  reg_psum_31_21;
assign out_psum_22 =  reg_psum_31_22;
assign out_psum_23 =  reg_psum_31_23;
assign out_psum_24 =  reg_psum_31_24;
assign out_psum_25 =  reg_psum_31_25;
assign out_psum_26 =  reg_psum_31_26;
assign out_psum_27 =  reg_psum_31_27;
assign out_psum_28 =  reg_psum_31_28;
assign out_psum_29 =  reg_psum_31_29;
assign out_psum_30 =  reg_psum_31_30;
assign out_psum_31 =  reg_psum_31_31;
wire signed[15:0]    fault_reg_psum_0_10;
wire signed[15:0]    fault_reg_psum_0_11;
wire signed[15:0]    fault_reg_psum_2_20;
wire signed[15:0]    fault_reg_psum_3_0;
wire signed[15:0]    fault_reg_psum_3_30;
wire signed[15:0]    fault_reg_psum_5_30;
wire signed[15:0]    fault_reg_psum_6_26;
wire signed[15:0]    fault_reg_psum_10_26;
wire signed[15:0]    fault_reg_psum_13_3;
wire signed[15:0]    fault_reg_psum_14_20;
wire signed[15:0]    fault_reg_psum_16_5;
wire signed[15:0]    fault_reg_psum_19_0;
wire signed[15:0]    fault_reg_psum_20_11;
wire signed[15:0]    fault_reg_psum_21_17;
wire signed[15:0]    fault_reg_psum_21_30;
wire signed[15:0]    fault_reg_psum_22_30;
wire signed[15:0]    fault_reg_psum_24_10;
wire signed[15:0]    fault_reg_psum_30_11;
assign fault_reg_psum_30_11 = reg_psum_30_11 | 16'b0000000001000000;
assign fault_reg_psum_24_10 = reg_psum_24_10 & 16'b1111111111110111;
assign fault_reg_psum_22_30 = reg_psum_22_30 | 16'b0000000000000001;
assign fault_reg_psum_21_30 = reg_psum_21_30 | 16'b0000000000000001;
assign fault_reg_psum_21_17 = reg_psum_21_17 & 16'b1111111111011111;
assign fault_reg_psum_20_11 = reg_psum_20_11 & 16'b1111111111011111;
assign fault_reg_psum_19_0 = reg_psum_19_0 | 16'b0000000000010000;
assign fault_reg_psum_16_5 = reg_psum_16_5 & 16'b1111110111111111;
assign fault_reg_psum_14_20 = reg_psum_14_20 & 16'b1111111101111111;
assign fault_reg_psum_13_3 = reg_psum_13_3 | 16'b0000000000000001;
assign fault_reg_psum_10_26 = reg_psum_10_26 & 16'b1111111011111111;
assign fault_reg_psum_6_26 = reg_psum_6_26 & 16'b1111101111111111;
assign fault_reg_psum_5_30 = reg_psum_5_30 | 16'b0000000001000000;
assign fault_reg_psum_3_0 = reg_psum_3_0 & 16'b1111111011111111;
assign fault_reg_psum_3_30 = reg_psum_3_30 | 16'b0000000000000010;
assign fault_reg_psum_2_20 = reg_psum_2_20 & 16'b1111111011111111;
assign fault_reg_psum_0_10 = reg_psum_0_10 | 16'b0000000000000100;
assign fault_reg_psum_0_11 = reg_psum_0_11 & 16'b1111111111111101;
PE U0_0( .activation_in(in_activation_0), .weight_in(in_weight_0), .partial_sum_in(in_psum_0), .reg_activation(reg_activation_0_0), .reg_weight(reg_weight_0_0), .reg_partial_sum(reg_psum_0_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_1( .activation_in(reg_activation_0_0), .weight_in(in_weight_1), .partial_sum_in(in_psum_1), .reg_activation(reg_activation_0_1), .reg_weight(reg_weight_0_1), .reg_partial_sum(reg_psum_0_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_2( .activation_in(reg_activation_0_1), .weight_in(in_weight_2), .partial_sum_in(in_psum_2), .reg_activation(reg_activation_0_2), .reg_weight(reg_weight_0_2), .reg_partial_sum(reg_psum_0_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_3( .activation_in(reg_activation_0_2), .weight_in(in_weight_3), .partial_sum_in(in_psum_3), .reg_activation(reg_activation_0_3), .reg_weight(reg_weight_0_3), .reg_partial_sum(reg_psum_0_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_4( .activation_in(reg_activation_0_3), .weight_in(in_weight_4), .partial_sum_in(in_psum_4), .reg_activation(reg_activation_0_4), .reg_weight(reg_weight_0_4), .reg_partial_sum(reg_psum_0_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_5( .activation_in(reg_activation_0_4), .weight_in(in_weight_5), .partial_sum_in(in_psum_5), .reg_activation(reg_activation_0_5), .reg_weight(reg_weight_0_5), .reg_partial_sum(reg_psum_0_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_6( .activation_in(reg_activation_0_5), .weight_in(in_weight_6), .partial_sum_in(in_psum_6), .reg_activation(reg_activation_0_6), .reg_weight(reg_weight_0_6), .reg_partial_sum(reg_psum_0_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_7( .activation_in(reg_activation_0_6), .weight_in(in_weight_7), .partial_sum_in(in_psum_7), .reg_activation(reg_activation_0_7), .reg_weight(reg_weight_0_7), .reg_partial_sum(reg_psum_0_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_8( .activation_in(reg_activation_0_7), .weight_in(in_weight_8), .partial_sum_in(in_psum_8), .reg_activation(reg_activation_0_8), .reg_weight(reg_weight_0_8), .reg_partial_sum(reg_psum_0_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_9( .activation_in(reg_activation_0_8), .weight_in(in_weight_9), .partial_sum_in(in_psum_9), .reg_activation(reg_activation_0_9), .reg_weight(reg_weight_0_9), .reg_partial_sum(reg_psum_0_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_10( .activation_in(reg_activation_0_9), .weight_in(in_weight_10), .partial_sum_in(in_psum_10), .reg_activation(reg_activation_0_10), .reg_weight(reg_weight_0_10), .reg_partial_sum(reg_psum_0_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_11( .activation_in(reg_activation_0_10), .weight_in(in_weight_11), .partial_sum_in(in_psum_11), .reg_activation(reg_activation_0_11), .reg_weight(reg_weight_0_11), .reg_partial_sum(reg_psum_0_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_12( .activation_in(reg_activation_0_11), .weight_in(in_weight_12), .partial_sum_in(in_psum_12), .reg_activation(reg_activation_0_12), .reg_weight(reg_weight_0_12), .reg_partial_sum(reg_psum_0_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_13( .activation_in(reg_activation_0_12), .weight_in(in_weight_13), .partial_sum_in(in_psum_13), .reg_activation(reg_activation_0_13), .reg_weight(reg_weight_0_13), .reg_partial_sum(reg_psum_0_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_14( .activation_in(reg_activation_0_13), .weight_in(in_weight_14), .partial_sum_in(in_psum_14), .reg_activation(reg_activation_0_14), .reg_weight(reg_weight_0_14), .reg_partial_sum(reg_psum_0_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_15( .activation_in(reg_activation_0_14), .weight_in(in_weight_15), .partial_sum_in(in_psum_15), .reg_activation(reg_activation_0_15), .reg_weight(reg_weight_0_15), .reg_partial_sum(reg_psum_0_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_16( .activation_in(reg_activation_0_15), .weight_in(in_weight_16), .partial_sum_in(in_psum_16), .reg_activation(reg_activation_0_16), .reg_weight(reg_weight_0_16), .reg_partial_sum(reg_psum_0_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_17( .activation_in(reg_activation_0_16), .weight_in(in_weight_17), .partial_sum_in(in_psum_17), .reg_activation(reg_activation_0_17), .reg_weight(reg_weight_0_17), .reg_partial_sum(reg_psum_0_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_18( .activation_in(reg_activation_0_17), .weight_in(in_weight_18), .partial_sum_in(in_psum_18), .reg_activation(reg_activation_0_18), .reg_weight(reg_weight_0_18), .reg_partial_sum(reg_psum_0_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_19( .activation_in(reg_activation_0_18), .weight_in(in_weight_19), .partial_sum_in(in_psum_19), .reg_activation(reg_activation_0_19), .reg_weight(reg_weight_0_19), .reg_partial_sum(reg_psum_0_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_20( .activation_in(reg_activation_0_19), .weight_in(in_weight_20), .partial_sum_in(in_psum_20), .reg_activation(reg_activation_0_20), .reg_weight(reg_weight_0_20), .reg_partial_sum(reg_psum_0_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_21( .activation_in(reg_activation_0_20), .weight_in(in_weight_21), .partial_sum_in(in_psum_21), .reg_activation(reg_activation_0_21), .reg_weight(reg_weight_0_21), .reg_partial_sum(reg_psum_0_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_22( .activation_in(reg_activation_0_21), .weight_in(in_weight_22), .partial_sum_in(in_psum_22), .reg_activation(reg_activation_0_22), .reg_weight(reg_weight_0_22), .reg_partial_sum(reg_psum_0_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_23( .activation_in(reg_activation_0_22), .weight_in(in_weight_23), .partial_sum_in(in_psum_23), .reg_activation(reg_activation_0_23), .reg_weight(reg_weight_0_23), .reg_partial_sum(reg_psum_0_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_24( .activation_in(reg_activation_0_23), .weight_in(in_weight_24), .partial_sum_in(in_psum_24), .reg_activation(reg_activation_0_24), .reg_weight(reg_weight_0_24), .reg_partial_sum(reg_psum_0_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_25( .activation_in(reg_activation_0_24), .weight_in(in_weight_25), .partial_sum_in(in_psum_25), .reg_activation(reg_activation_0_25), .reg_weight(reg_weight_0_25), .reg_partial_sum(reg_psum_0_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_26( .activation_in(reg_activation_0_25), .weight_in(in_weight_26), .partial_sum_in(in_psum_26), .reg_activation(reg_activation_0_26), .reg_weight(reg_weight_0_26), .reg_partial_sum(reg_psum_0_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_27( .activation_in(reg_activation_0_26), .weight_in(in_weight_27), .partial_sum_in(in_psum_27), .reg_activation(reg_activation_0_27), .reg_weight(reg_weight_0_27), .reg_partial_sum(reg_psum_0_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_28( .activation_in(reg_activation_0_27), .weight_in(in_weight_28), .partial_sum_in(in_psum_28), .reg_activation(reg_activation_0_28), .reg_weight(reg_weight_0_28), .reg_partial_sum(reg_psum_0_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_29( .activation_in(reg_activation_0_28), .weight_in(in_weight_29), .partial_sum_in(in_psum_29), .reg_activation(reg_activation_0_29), .reg_weight(reg_weight_0_29), .reg_partial_sum(reg_psum_0_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_30( .activation_in(reg_activation_0_29), .weight_in(in_weight_30), .partial_sum_in(in_psum_30), .reg_activation(reg_activation_0_30), .reg_weight(reg_weight_0_30), .reg_partial_sum(reg_psum_0_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U0_31( .activation_in(reg_activation_0_30), .weight_in(in_weight_31), .partial_sum_in(in_psum_31), .reg_weight(reg_weight_0_31), .reg_partial_sum(reg_psum_0_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_0( .activation_in(in_activation_1), .weight_in(reg_weight_0_0), .partial_sum_in(reg_psum_0_0), .reg_activation(reg_activation_1_0), .reg_weight(reg_weight_1_0), .reg_partial_sum(reg_psum_1_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_1( .activation_in(reg_activation_1_0), .weight_in(reg_weight_0_1), .partial_sum_in(reg_psum_0_1), .reg_activation(reg_activation_1_1), .reg_weight(reg_weight_1_1), .reg_partial_sum(reg_psum_1_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_2( .activation_in(reg_activation_1_1), .weight_in(reg_weight_0_2), .partial_sum_in(reg_psum_0_2), .reg_activation(reg_activation_1_2), .reg_weight(reg_weight_1_2), .reg_partial_sum(reg_psum_1_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_3( .activation_in(reg_activation_1_2), .weight_in(reg_weight_0_3), .partial_sum_in(reg_psum_0_3), .reg_activation(reg_activation_1_3), .reg_weight(reg_weight_1_3), .reg_partial_sum(reg_psum_1_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_4( .activation_in(reg_activation_1_3), .weight_in(reg_weight_0_4), .partial_sum_in(reg_psum_0_4), .reg_activation(reg_activation_1_4), .reg_weight(reg_weight_1_4), .reg_partial_sum(reg_psum_1_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_5( .activation_in(reg_activation_1_4), .weight_in(reg_weight_0_5), .partial_sum_in(reg_psum_0_5), .reg_activation(reg_activation_1_5), .reg_weight(reg_weight_1_5), .reg_partial_sum(reg_psum_1_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_6( .activation_in(reg_activation_1_5), .weight_in(reg_weight_0_6), .partial_sum_in(reg_psum_0_6), .reg_activation(reg_activation_1_6), .reg_weight(reg_weight_1_6), .reg_partial_sum(reg_psum_1_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_7( .activation_in(reg_activation_1_6), .weight_in(reg_weight_0_7), .partial_sum_in(reg_psum_0_7), .reg_activation(reg_activation_1_7), .reg_weight(reg_weight_1_7), .reg_partial_sum(reg_psum_1_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_8( .activation_in(reg_activation_1_7), .weight_in(reg_weight_0_8), .partial_sum_in(reg_psum_0_8), .reg_activation(reg_activation_1_8), .reg_weight(reg_weight_1_8), .reg_partial_sum(reg_psum_1_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_9( .activation_in(reg_activation_1_8), .weight_in(reg_weight_0_9), .partial_sum_in(reg_psum_0_9), .reg_activation(reg_activation_1_9), .reg_weight(reg_weight_1_9), .reg_partial_sum(reg_psum_1_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_10( .activation_in(reg_activation_1_9), .weight_in(reg_weight_0_10), .partial_sum_in(fault_reg_psum_0_10), .reg_activation(reg_activation_1_10), .reg_weight(reg_weight_1_10), .reg_partial_sum(reg_psum_1_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_11( .activation_in(reg_activation_1_10), .weight_in(reg_weight_0_11), .partial_sum_in(fault_reg_psum_0_11), .reg_activation(reg_activation_1_11), .reg_weight(reg_weight_1_11), .reg_partial_sum(reg_psum_1_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_12( .activation_in(reg_activation_1_11), .weight_in(reg_weight_0_12), .partial_sum_in(reg_psum_0_12), .reg_activation(reg_activation_1_12), .reg_weight(reg_weight_1_12), .reg_partial_sum(reg_psum_1_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_13( .activation_in(reg_activation_1_12), .weight_in(reg_weight_0_13), .partial_sum_in(reg_psum_0_13), .reg_activation(reg_activation_1_13), .reg_weight(reg_weight_1_13), .reg_partial_sum(reg_psum_1_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_14( .activation_in(reg_activation_1_13), .weight_in(reg_weight_0_14), .partial_sum_in(reg_psum_0_14), .reg_activation(reg_activation_1_14), .reg_weight(reg_weight_1_14), .reg_partial_sum(reg_psum_1_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_15( .activation_in(reg_activation_1_14), .weight_in(reg_weight_0_15), .partial_sum_in(reg_psum_0_15), .reg_activation(reg_activation_1_15), .reg_weight(reg_weight_1_15), .reg_partial_sum(reg_psum_1_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_16( .activation_in(reg_activation_1_15), .weight_in(reg_weight_0_16), .partial_sum_in(reg_psum_0_16), .reg_activation(reg_activation_1_16), .reg_weight(reg_weight_1_16), .reg_partial_sum(reg_psum_1_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_17( .activation_in(reg_activation_1_16), .weight_in(reg_weight_0_17), .partial_sum_in(reg_psum_0_17), .reg_activation(reg_activation_1_17), .reg_weight(reg_weight_1_17), .reg_partial_sum(reg_psum_1_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_18( .activation_in(reg_activation_1_17), .weight_in(reg_weight_0_18), .partial_sum_in(reg_psum_0_18), .reg_activation(reg_activation_1_18), .reg_weight(reg_weight_1_18), .reg_partial_sum(reg_psum_1_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_19( .activation_in(reg_activation_1_18), .weight_in(reg_weight_0_19), .partial_sum_in(reg_psum_0_19), .reg_activation(reg_activation_1_19), .reg_weight(reg_weight_1_19), .reg_partial_sum(reg_psum_1_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_20( .activation_in(reg_activation_1_19), .weight_in(reg_weight_0_20), .partial_sum_in(reg_psum_0_20), .reg_activation(reg_activation_1_20), .reg_weight(reg_weight_1_20), .reg_partial_sum(reg_psum_1_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_21( .activation_in(reg_activation_1_20), .weight_in(reg_weight_0_21), .partial_sum_in(reg_psum_0_21), .reg_activation(reg_activation_1_21), .reg_weight(reg_weight_1_21), .reg_partial_sum(reg_psum_1_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_22( .activation_in(reg_activation_1_21), .weight_in(reg_weight_0_22), .partial_sum_in(reg_psum_0_22), .reg_activation(reg_activation_1_22), .reg_weight(reg_weight_1_22), .reg_partial_sum(reg_psum_1_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_23( .activation_in(reg_activation_1_22), .weight_in(reg_weight_0_23), .partial_sum_in(reg_psum_0_23), .reg_activation(reg_activation_1_23), .reg_weight(reg_weight_1_23), .reg_partial_sum(reg_psum_1_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_24( .activation_in(reg_activation_1_23), .weight_in(reg_weight_0_24), .partial_sum_in(reg_psum_0_24), .reg_activation(reg_activation_1_24), .reg_weight(reg_weight_1_24), .reg_partial_sum(reg_psum_1_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_25( .activation_in(reg_activation_1_24), .weight_in(reg_weight_0_25), .partial_sum_in(reg_psum_0_25), .reg_activation(reg_activation_1_25), .reg_weight(reg_weight_1_25), .reg_partial_sum(reg_psum_1_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_26( .activation_in(reg_activation_1_25), .weight_in(reg_weight_0_26), .partial_sum_in(reg_psum_0_26), .reg_activation(reg_activation_1_26), .reg_weight(reg_weight_1_26), .reg_partial_sum(reg_psum_1_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_27( .activation_in(reg_activation_1_26), .weight_in(reg_weight_0_27), .partial_sum_in(reg_psum_0_27), .reg_activation(reg_activation_1_27), .reg_weight(reg_weight_1_27), .reg_partial_sum(reg_psum_1_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_28( .activation_in(reg_activation_1_27), .weight_in(reg_weight_0_28), .partial_sum_in(reg_psum_0_28), .reg_activation(reg_activation_1_28), .reg_weight(reg_weight_1_28), .reg_partial_sum(reg_psum_1_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_29( .activation_in(reg_activation_1_28), .weight_in(reg_weight_0_29), .partial_sum_in(reg_psum_0_29), .reg_activation(reg_activation_1_29), .reg_weight(reg_weight_1_29), .reg_partial_sum(reg_psum_1_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_30( .activation_in(reg_activation_1_29), .weight_in(reg_weight_0_30), .partial_sum_in(reg_psum_0_30), .reg_activation(reg_activation_1_30), .reg_weight(reg_weight_1_30), .reg_partial_sum(reg_psum_1_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U1_31( .activation_in(reg_activation_1_30), .weight_in(reg_weight_0_31), .partial_sum_in(reg_psum_0_31), .reg_weight(reg_weight_1_31), .reg_partial_sum(reg_psum_1_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_0( .activation_in(in_activation_2), .weight_in(reg_weight_1_0), .partial_sum_in(reg_psum_1_0), .reg_activation(reg_activation_2_0), .reg_weight(reg_weight_2_0), .reg_partial_sum(reg_psum_2_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_1( .activation_in(reg_activation_2_0), .weight_in(reg_weight_1_1), .partial_sum_in(reg_psum_1_1), .reg_activation(reg_activation_2_1), .reg_weight(reg_weight_2_1), .reg_partial_sum(reg_psum_2_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_2( .activation_in(reg_activation_2_1), .weight_in(reg_weight_1_2), .partial_sum_in(reg_psum_1_2), .reg_activation(reg_activation_2_2), .reg_weight(reg_weight_2_2), .reg_partial_sum(reg_psum_2_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_3( .activation_in(reg_activation_2_2), .weight_in(reg_weight_1_3), .partial_sum_in(reg_psum_1_3), .reg_activation(reg_activation_2_3), .reg_weight(reg_weight_2_3), .reg_partial_sum(reg_psum_2_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_4( .activation_in(reg_activation_2_3), .weight_in(reg_weight_1_4), .partial_sum_in(reg_psum_1_4), .reg_activation(reg_activation_2_4), .reg_weight(reg_weight_2_4), .reg_partial_sum(reg_psum_2_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_5( .activation_in(reg_activation_2_4), .weight_in(reg_weight_1_5), .partial_sum_in(reg_psum_1_5), .reg_activation(reg_activation_2_5), .reg_weight(reg_weight_2_5), .reg_partial_sum(reg_psum_2_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_6( .activation_in(reg_activation_2_5), .weight_in(reg_weight_1_6), .partial_sum_in(reg_psum_1_6), .reg_activation(reg_activation_2_6), .reg_weight(reg_weight_2_6), .reg_partial_sum(reg_psum_2_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_7( .activation_in(reg_activation_2_6), .weight_in(reg_weight_1_7), .partial_sum_in(reg_psum_1_7), .reg_activation(reg_activation_2_7), .reg_weight(reg_weight_2_7), .reg_partial_sum(reg_psum_2_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_8( .activation_in(reg_activation_2_7), .weight_in(reg_weight_1_8), .partial_sum_in(reg_psum_1_8), .reg_activation(reg_activation_2_8), .reg_weight(reg_weight_2_8), .reg_partial_sum(reg_psum_2_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_9( .activation_in(reg_activation_2_8), .weight_in(reg_weight_1_9), .partial_sum_in(reg_psum_1_9), .reg_activation(reg_activation_2_9), .reg_weight(reg_weight_2_9), .reg_partial_sum(reg_psum_2_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_10( .activation_in(reg_activation_2_9), .weight_in(reg_weight_1_10), .partial_sum_in(reg_psum_1_10), .reg_activation(reg_activation_2_10), .reg_weight(reg_weight_2_10), .reg_partial_sum(reg_psum_2_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_11( .activation_in(reg_activation_2_10), .weight_in(reg_weight_1_11), .partial_sum_in(reg_psum_1_11), .reg_activation(reg_activation_2_11), .reg_weight(reg_weight_2_11), .reg_partial_sum(reg_psum_2_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_12( .activation_in(reg_activation_2_11), .weight_in(reg_weight_1_12), .partial_sum_in(reg_psum_1_12), .reg_activation(reg_activation_2_12), .reg_weight(reg_weight_2_12), .reg_partial_sum(reg_psum_2_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_13( .activation_in(reg_activation_2_12), .weight_in(reg_weight_1_13), .partial_sum_in(reg_psum_1_13), .reg_activation(reg_activation_2_13), .reg_weight(reg_weight_2_13), .reg_partial_sum(reg_psum_2_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_14( .activation_in(reg_activation_2_13), .weight_in(reg_weight_1_14), .partial_sum_in(reg_psum_1_14), .reg_activation(reg_activation_2_14), .reg_weight(reg_weight_2_14), .reg_partial_sum(reg_psum_2_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_15( .activation_in(reg_activation_2_14), .weight_in(reg_weight_1_15), .partial_sum_in(reg_psum_1_15), .reg_activation(reg_activation_2_15), .reg_weight(reg_weight_2_15), .reg_partial_sum(reg_psum_2_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_16( .activation_in(reg_activation_2_15), .weight_in(reg_weight_1_16), .partial_sum_in(reg_psum_1_16), .reg_activation(reg_activation_2_16), .reg_weight(reg_weight_2_16), .reg_partial_sum(reg_psum_2_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_17( .activation_in(reg_activation_2_16), .weight_in(reg_weight_1_17), .partial_sum_in(reg_psum_1_17), .reg_activation(reg_activation_2_17), .reg_weight(reg_weight_2_17), .reg_partial_sum(reg_psum_2_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_18( .activation_in(reg_activation_2_17), .weight_in(reg_weight_1_18), .partial_sum_in(reg_psum_1_18), .reg_activation(reg_activation_2_18), .reg_weight(reg_weight_2_18), .reg_partial_sum(reg_psum_2_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_19( .activation_in(reg_activation_2_18), .weight_in(reg_weight_1_19), .partial_sum_in(reg_psum_1_19), .reg_activation(reg_activation_2_19), .reg_weight(reg_weight_2_19), .reg_partial_sum(reg_psum_2_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_20( .activation_in(reg_activation_2_19), .weight_in(reg_weight_1_20), .partial_sum_in(reg_psum_1_20), .reg_activation(reg_activation_2_20), .reg_weight(reg_weight_2_20), .reg_partial_sum(reg_psum_2_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_21( .activation_in(reg_activation_2_20), .weight_in(reg_weight_1_21), .partial_sum_in(reg_psum_1_21), .reg_activation(reg_activation_2_21), .reg_weight(reg_weight_2_21), .reg_partial_sum(reg_psum_2_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_22( .activation_in(reg_activation_2_21), .weight_in(reg_weight_1_22), .partial_sum_in(reg_psum_1_22), .reg_activation(reg_activation_2_22), .reg_weight(reg_weight_2_22), .reg_partial_sum(reg_psum_2_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_23( .activation_in(reg_activation_2_22), .weight_in(reg_weight_1_23), .partial_sum_in(reg_psum_1_23), .reg_activation(reg_activation_2_23), .reg_weight(reg_weight_2_23), .reg_partial_sum(reg_psum_2_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_24( .activation_in(reg_activation_2_23), .weight_in(reg_weight_1_24), .partial_sum_in(reg_psum_1_24), .reg_activation(reg_activation_2_24), .reg_weight(reg_weight_2_24), .reg_partial_sum(reg_psum_2_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_25( .activation_in(reg_activation_2_24), .weight_in(reg_weight_1_25), .partial_sum_in(reg_psum_1_25), .reg_activation(reg_activation_2_25), .reg_weight(reg_weight_2_25), .reg_partial_sum(reg_psum_2_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_26( .activation_in(reg_activation_2_25), .weight_in(reg_weight_1_26), .partial_sum_in(reg_psum_1_26), .reg_activation(reg_activation_2_26), .reg_weight(reg_weight_2_26), .reg_partial_sum(reg_psum_2_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_27( .activation_in(reg_activation_2_26), .weight_in(reg_weight_1_27), .partial_sum_in(reg_psum_1_27), .reg_activation(reg_activation_2_27), .reg_weight(reg_weight_2_27), .reg_partial_sum(reg_psum_2_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_28( .activation_in(reg_activation_2_27), .weight_in(reg_weight_1_28), .partial_sum_in(reg_psum_1_28), .reg_activation(reg_activation_2_28), .reg_weight(reg_weight_2_28), .reg_partial_sum(reg_psum_2_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_29( .activation_in(reg_activation_2_28), .weight_in(reg_weight_1_29), .partial_sum_in(reg_psum_1_29), .reg_activation(reg_activation_2_29), .reg_weight(reg_weight_2_29), .reg_partial_sum(reg_psum_2_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_30( .activation_in(reg_activation_2_29), .weight_in(reg_weight_1_30), .partial_sum_in(reg_psum_1_30), .reg_activation(reg_activation_2_30), .reg_weight(reg_weight_2_30), .reg_partial_sum(reg_psum_2_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U2_31( .activation_in(reg_activation_2_30), .weight_in(reg_weight_1_31), .partial_sum_in(reg_psum_1_31), .reg_weight(reg_weight_2_31), .reg_partial_sum(reg_psum_2_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_0( .activation_in(in_activation_3), .weight_in(reg_weight_2_0), .partial_sum_in(reg_psum_2_0), .reg_activation(reg_activation_3_0), .reg_weight(reg_weight_3_0), .reg_partial_sum(reg_psum_3_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_1( .activation_in(reg_activation_3_0), .weight_in(reg_weight_2_1), .partial_sum_in(reg_psum_2_1), .reg_activation(reg_activation_3_1), .reg_weight(reg_weight_3_1), .reg_partial_sum(reg_psum_3_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_2( .activation_in(reg_activation_3_1), .weight_in(reg_weight_2_2), .partial_sum_in(reg_psum_2_2), .reg_activation(reg_activation_3_2), .reg_weight(reg_weight_3_2), .reg_partial_sum(reg_psum_3_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_3( .activation_in(reg_activation_3_2), .weight_in(reg_weight_2_3), .partial_sum_in(reg_psum_2_3), .reg_activation(reg_activation_3_3), .reg_weight(reg_weight_3_3), .reg_partial_sum(reg_psum_3_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_4( .activation_in(reg_activation_3_3), .weight_in(reg_weight_2_4), .partial_sum_in(reg_psum_2_4), .reg_activation(reg_activation_3_4), .reg_weight(reg_weight_3_4), .reg_partial_sum(reg_psum_3_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_5( .activation_in(reg_activation_3_4), .weight_in(reg_weight_2_5), .partial_sum_in(reg_psum_2_5), .reg_activation(reg_activation_3_5), .reg_weight(reg_weight_3_5), .reg_partial_sum(reg_psum_3_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_6( .activation_in(reg_activation_3_5), .weight_in(reg_weight_2_6), .partial_sum_in(reg_psum_2_6), .reg_activation(reg_activation_3_6), .reg_weight(reg_weight_3_6), .reg_partial_sum(reg_psum_3_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_7( .activation_in(reg_activation_3_6), .weight_in(reg_weight_2_7), .partial_sum_in(reg_psum_2_7), .reg_activation(reg_activation_3_7), .reg_weight(reg_weight_3_7), .reg_partial_sum(reg_psum_3_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_8( .activation_in(reg_activation_3_7), .weight_in(reg_weight_2_8), .partial_sum_in(reg_psum_2_8), .reg_activation(reg_activation_3_8), .reg_weight(reg_weight_3_8), .reg_partial_sum(reg_psum_3_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_9( .activation_in(reg_activation_3_8), .weight_in(reg_weight_2_9), .partial_sum_in(reg_psum_2_9), .reg_activation(reg_activation_3_9), .reg_weight(reg_weight_3_9), .reg_partial_sum(reg_psum_3_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_10( .activation_in(reg_activation_3_9), .weight_in(reg_weight_2_10), .partial_sum_in(reg_psum_2_10), .reg_activation(reg_activation_3_10), .reg_weight(reg_weight_3_10), .reg_partial_sum(reg_psum_3_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_11( .activation_in(reg_activation_3_10), .weight_in(reg_weight_2_11), .partial_sum_in(reg_psum_2_11), .reg_activation(reg_activation_3_11), .reg_weight(reg_weight_3_11), .reg_partial_sum(reg_psum_3_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_12( .activation_in(reg_activation_3_11), .weight_in(reg_weight_2_12), .partial_sum_in(reg_psum_2_12), .reg_activation(reg_activation_3_12), .reg_weight(reg_weight_3_12), .reg_partial_sum(reg_psum_3_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_13( .activation_in(reg_activation_3_12), .weight_in(reg_weight_2_13), .partial_sum_in(reg_psum_2_13), .reg_activation(reg_activation_3_13), .reg_weight(reg_weight_3_13), .reg_partial_sum(reg_psum_3_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_14( .activation_in(reg_activation_3_13), .weight_in(reg_weight_2_14), .partial_sum_in(reg_psum_2_14), .reg_activation(reg_activation_3_14), .reg_weight(reg_weight_3_14), .reg_partial_sum(reg_psum_3_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_15( .activation_in(reg_activation_3_14), .weight_in(reg_weight_2_15), .partial_sum_in(reg_psum_2_15), .reg_activation(reg_activation_3_15), .reg_weight(reg_weight_3_15), .reg_partial_sum(reg_psum_3_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_16( .activation_in(reg_activation_3_15), .weight_in(reg_weight_2_16), .partial_sum_in(reg_psum_2_16), .reg_activation(reg_activation_3_16), .reg_weight(reg_weight_3_16), .reg_partial_sum(reg_psum_3_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_17( .activation_in(reg_activation_3_16), .weight_in(reg_weight_2_17), .partial_sum_in(reg_psum_2_17), .reg_activation(reg_activation_3_17), .reg_weight(reg_weight_3_17), .reg_partial_sum(reg_psum_3_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_18( .activation_in(reg_activation_3_17), .weight_in(reg_weight_2_18), .partial_sum_in(reg_psum_2_18), .reg_activation(reg_activation_3_18), .reg_weight(reg_weight_3_18), .reg_partial_sum(reg_psum_3_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_19( .activation_in(reg_activation_3_18), .weight_in(reg_weight_2_19), .partial_sum_in(reg_psum_2_19), .reg_activation(reg_activation_3_19), .reg_weight(reg_weight_3_19), .reg_partial_sum(reg_psum_3_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_20( .activation_in(reg_activation_3_19), .weight_in(reg_weight_2_20), .partial_sum_in(fault_reg_psum_2_20), .reg_activation(reg_activation_3_20), .reg_weight(reg_weight_3_20), .reg_partial_sum(reg_psum_3_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_21( .activation_in(reg_activation_3_20), .weight_in(reg_weight_2_21), .partial_sum_in(reg_psum_2_21), .reg_activation(reg_activation_3_21), .reg_weight(reg_weight_3_21), .reg_partial_sum(reg_psum_3_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_22( .activation_in(reg_activation_3_21), .weight_in(reg_weight_2_22), .partial_sum_in(reg_psum_2_22), .reg_activation(reg_activation_3_22), .reg_weight(reg_weight_3_22), .reg_partial_sum(reg_psum_3_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_23( .activation_in(reg_activation_3_22), .weight_in(reg_weight_2_23), .partial_sum_in(reg_psum_2_23), .reg_activation(reg_activation_3_23), .reg_weight(reg_weight_3_23), .reg_partial_sum(reg_psum_3_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_24( .activation_in(reg_activation_3_23), .weight_in(reg_weight_2_24), .partial_sum_in(reg_psum_2_24), .reg_activation(reg_activation_3_24), .reg_weight(reg_weight_3_24), .reg_partial_sum(reg_psum_3_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_25( .activation_in(reg_activation_3_24), .weight_in(reg_weight_2_25), .partial_sum_in(reg_psum_2_25), .reg_activation(reg_activation_3_25), .reg_weight(reg_weight_3_25), .reg_partial_sum(reg_psum_3_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_26( .activation_in(reg_activation_3_25), .weight_in(reg_weight_2_26), .partial_sum_in(reg_psum_2_26), .reg_activation(reg_activation_3_26), .reg_weight(reg_weight_3_26), .reg_partial_sum(reg_psum_3_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_27( .activation_in(reg_activation_3_26), .weight_in(reg_weight_2_27), .partial_sum_in(reg_psum_2_27), .reg_activation(reg_activation_3_27), .reg_weight(reg_weight_3_27), .reg_partial_sum(reg_psum_3_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_28( .activation_in(reg_activation_3_27), .weight_in(reg_weight_2_28), .partial_sum_in(reg_psum_2_28), .reg_activation(reg_activation_3_28), .reg_weight(reg_weight_3_28), .reg_partial_sum(reg_psum_3_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_29( .activation_in(reg_activation_3_28), .weight_in(reg_weight_2_29), .partial_sum_in(reg_psum_2_29), .reg_activation(reg_activation_3_29), .reg_weight(reg_weight_3_29), .reg_partial_sum(reg_psum_3_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_30( .activation_in(reg_activation_3_29), .weight_in(reg_weight_2_30), .partial_sum_in(reg_psum_2_30), .reg_activation(reg_activation_3_30), .reg_weight(reg_weight_3_30), .reg_partial_sum(reg_psum_3_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U3_31( .activation_in(reg_activation_3_30), .weight_in(reg_weight_2_31), .partial_sum_in(reg_psum_2_31), .reg_weight(reg_weight_3_31), .reg_partial_sum(reg_psum_3_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_0( .activation_in(in_activation_4), .weight_in(reg_weight_3_0), .partial_sum_in(fault_reg_psum_3_0), .reg_activation(reg_activation_4_0), .reg_weight(reg_weight_4_0), .reg_partial_sum(reg_psum_4_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_1( .activation_in(reg_activation_4_0), .weight_in(reg_weight_3_1), .partial_sum_in(reg_psum_3_1), .reg_activation(reg_activation_4_1), .reg_weight(reg_weight_4_1), .reg_partial_sum(reg_psum_4_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_2( .activation_in(reg_activation_4_1), .weight_in(reg_weight_3_2), .partial_sum_in(reg_psum_3_2), .reg_activation(reg_activation_4_2), .reg_weight(reg_weight_4_2), .reg_partial_sum(reg_psum_4_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_3( .activation_in(reg_activation_4_2), .weight_in(reg_weight_3_3), .partial_sum_in(reg_psum_3_3), .reg_activation(reg_activation_4_3), .reg_weight(reg_weight_4_3), .reg_partial_sum(reg_psum_4_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_4( .activation_in(reg_activation_4_3), .weight_in(reg_weight_3_4), .partial_sum_in(reg_psum_3_4), .reg_activation(reg_activation_4_4), .reg_weight(reg_weight_4_4), .reg_partial_sum(reg_psum_4_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_5( .activation_in(reg_activation_4_4), .weight_in(reg_weight_3_5), .partial_sum_in(reg_psum_3_5), .reg_activation(reg_activation_4_5), .reg_weight(reg_weight_4_5), .reg_partial_sum(reg_psum_4_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_6( .activation_in(reg_activation_4_5), .weight_in(reg_weight_3_6), .partial_sum_in(reg_psum_3_6), .reg_activation(reg_activation_4_6), .reg_weight(reg_weight_4_6), .reg_partial_sum(reg_psum_4_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_7( .activation_in(reg_activation_4_6), .weight_in(reg_weight_3_7), .partial_sum_in(reg_psum_3_7), .reg_activation(reg_activation_4_7), .reg_weight(reg_weight_4_7), .reg_partial_sum(reg_psum_4_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_8( .activation_in(reg_activation_4_7), .weight_in(reg_weight_3_8), .partial_sum_in(reg_psum_3_8), .reg_activation(reg_activation_4_8), .reg_weight(reg_weight_4_8), .reg_partial_sum(reg_psum_4_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_9( .activation_in(reg_activation_4_8), .weight_in(reg_weight_3_9), .partial_sum_in(reg_psum_3_9), .reg_activation(reg_activation_4_9), .reg_weight(reg_weight_4_9), .reg_partial_sum(reg_psum_4_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_10( .activation_in(reg_activation_4_9), .weight_in(reg_weight_3_10), .partial_sum_in(reg_psum_3_10), .reg_activation(reg_activation_4_10), .reg_weight(reg_weight_4_10), .reg_partial_sum(reg_psum_4_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_11( .activation_in(reg_activation_4_10), .weight_in(reg_weight_3_11), .partial_sum_in(reg_psum_3_11), .reg_activation(reg_activation_4_11), .reg_weight(reg_weight_4_11), .reg_partial_sum(reg_psum_4_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_12( .activation_in(reg_activation_4_11), .weight_in(reg_weight_3_12), .partial_sum_in(reg_psum_3_12), .reg_activation(reg_activation_4_12), .reg_weight(reg_weight_4_12), .reg_partial_sum(reg_psum_4_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_13( .activation_in(reg_activation_4_12), .weight_in(reg_weight_3_13), .partial_sum_in(reg_psum_3_13), .reg_activation(reg_activation_4_13), .reg_weight(reg_weight_4_13), .reg_partial_sum(reg_psum_4_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_14( .activation_in(reg_activation_4_13), .weight_in(reg_weight_3_14), .partial_sum_in(reg_psum_3_14), .reg_activation(reg_activation_4_14), .reg_weight(reg_weight_4_14), .reg_partial_sum(reg_psum_4_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_15( .activation_in(reg_activation_4_14), .weight_in(reg_weight_3_15), .partial_sum_in(reg_psum_3_15), .reg_activation(reg_activation_4_15), .reg_weight(reg_weight_4_15), .reg_partial_sum(reg_psum_4_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_16( .activation_in(reg_activation_4_15), .weight_in(reg_weight_3_16), .partial_sum_in(reg_psum_3_16), .reg_activation(reg_activation_4_16), .reg_weight(reg_weight_4_16), .reg_partial_sum(reg_psum_4_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_17( .activation_in(reg_activation_4_16), .weight_in(reg_weight_3_17), .partial_sum_in(reg_psum_3_17), .reg_activation(reg_activation_4_17), .reg_weight(reg_weight_4_17), .reg_partial_sum(reg_psum_4_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_18( .activation_in(reg_activation_4_17), .weight_in(reg_weight_3_18), .partial_sum_in(reg_psum_3_18), .reg_activation(reg_activation_4_18), .reg_weight(reg_weight_4_18), .reg_partial_sum(reg_psum_4_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_19( .activation_in(reg_activation_4_18), .weight_in(reg_weight_3_19), .partial_sum_in(reg_psum_3_19), .reg_activation(reg_activation_4_19), .reg_weight(reg_weight_4_19), .reg_partial_sum(reg_psum_4_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_20( .activation_in(reg_activation_4_19), .weight_in(reg_weight_3_20), .partial_sum_in(reg_psum_3_20), .reg_activation(reg_activation_4_20), .reg_weight(reg_weight_4_20), .reg_partial_sum(reg_psum_4_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_21( .activation_in(reg_activation_4_20), .weight_in(reg_weight_3_21), .partial_sum_in(reg_psum_3_21), .reg_activation(reg_activation_4_21), .reg_weight(reg_weight_4_21), .reg_partial_sum(reg_psum_4_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_22( .activation_in(reg_activation_4_21), .weight_in(reg_weight_3_22), .partial_sum_in(reg_psum_3_22), .reg_activation(reg_activation_4_22), .reg_weight(reg_weight_4_22), .reg_partial_sum(reg_psum_4_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_23( .activation_in(reg_activation_4_22), .weight_in(reg_weight_3_23), .partial_sum_in(reg_psum_3_23), .reg_activation(reg_activation_4_23), .reg_weight(reg_weight_4_23), .reg_partial_sum(reg_psum_4_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_24( .activation_in(reg_activation_4_23), .weight_in(reg_weight_3_24), .partial_sum_in(reg_psum_3_24), .reg_activation(reg_activation_4_24), .reg_weight(reg_weight_4_24), .reg_partial_sum(reg_psum_4_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_25( .activation_in(reg_activation_4_24), .weight_in(reg_weight_3_25), .partial_sum_in(reg_psum_3_25), .reg_activation(reg_activation_4_25), .reg_weight(reg_weight_4_25), .reg_partial_sum(reg_psum_4_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_26( .activation_in(reg_activation_4_25), .weight_in(reg_weight_3_26), .partial_sum_in(reg_psum_3_26), .reg_activation(reg_activation_4_26), .reg_weight(reg_weight_4_26), .reg_partial_sum(reg_psum_4_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_27( .activation_in(reg_activation_4_26), .weight_in(reg_weight_3_27), .partial_sum_in(reg_psum_3_27), .reg_activation(reg_activation_4_27), .reg_weight(reg_weight_4_27), .reg_partial_sum(reg_psum_4_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_28( .activation_in(reg_activation_4_27), .weight_in(reg_weight_3_28), .partial_sum_in(reg_psum_3_28), .reg_activation(reg_activation_4_28), .reg_weight(reg_weight_4_28), .reg_partial_sum(reg_psum_4_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_29( .activation_in(reg_activation_4_28), .weight_in(reg_weight_3_29), .partial_sum_in(reg_psum_3_29), .reg_activation(reg_activation_4_29), .reg_weight(reg_weight_4_29), .reg_partial_sum(reg_psum_4_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_30( .activation_in(reg_activation_4_29), .weight_in(reg_weight_3_30), .partial_sum_in(fault_reg_psum_3_30), .reg_activation(reg_activation_4_30), .reg_weight(reg_weight_4_30), .reg_partial_sum(reg_psum_4_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U4_31( .activation_in(reg_activation_4_30), .weight_in(reg_weight_3_31), .partial_sum_in(reg_psum_3_31), .reg_weight(reg_weight_4_31), .reg_partial_sum(reg_psum_4_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_0( .activation_in(in_activation_5), .weight_in(reg_weight_4_0), .partial_sum_in(reg_psum_4_0), .reg_activation(reg_activation_5_0), .reg_weight(reg_weight_5_0), .reg_partial_sum(reg_psum_5_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_1( .activation_in(reg_activation_5_0), .weight_in(reg_weight_4_1), .partial_sum_in(reg_psum_4_1), .reg_activation(reg_activation_5_1), .reg_weight(reg_weight_5_1), .reg_partial_sum(reg_psum_5_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_2( .activation_in(reg_activation_5_1), .weight_in(reg_weight_4_2), .partial_sum_in(reg_psum_4_2), .reg_activation(reg_activation_5_2), .reg_weight(reg_weight_5_2), .reg_partial_sum(reg_psum_5_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_3( .activation_in(reg_activation_5_2), .weight_in(reg_weight_4_3), .partial_sum_in(reg_psum_4_3), .reg_activation(reg_activation_5_3), .reg_weight(reg_weight_5_3), .reg_partial_sum(reg_psum_5_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_4( .activation_in(reg_activation_5_3), .weight_in(reg_weight_4_4), .partial_sum_in(reg_psum_4_4), .reg_activation(reg_activation_5_4), .reg_weight(reg_weight_5_4), .reg_partial_sum(reg_psum_5_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_5( .activation_in(reg_activation_5_4), .weight_in(reg_weight_4_5), .partial_sum_in(reg_psum_4_5), .reg_activation(reg_activation_5_5), .reg_weight(reg_weight_5_5), .reg_partial_sum(reg_psum_5_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_6( .activation_in(reg_activation_5_5), .weight_in(reg_weight_4_6), .partial_sum_in(reg_psum_4_6), .reg_activation(reg_activation_5_6), .reg_weight(reg_weight_5_6), .reg_partial_sum(reg_psum_5_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_7( .activation_in(reg_activation_5_6), .weight_in(reg_weight_4_7), .partial_sum_in(reg_psum_4_7), .reg_activation(reg_activation_5_7), .reg_weight(reg_weight_5_7), .reg_partial_sum(reg_psum_5_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_8( .activation_in(reg_activation_5_7), .weight_in(reg_weight_4_8), .partial_sum_in(reg_psum_4_8), .reg_activation(reg_activation_5_8), .reg_weight(reg_weight_5_8), .reg_partial_sum(reg_psum_5_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_9( .activation_in(reg_activation_5_8), .weight_in(reg_weight_4_9), .partial_sum_in(reg_psum_4_9), .reg_activation(reg_activation_5_9), .reg_weight(reg_weight_5_9), .reg_partial_sum(reg_psum_5_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_10( .activation_in(reg_activation_5_9), .weight_in(reg_weight_4_10), .partial_sum_in(reg_psum_4_10), .reg_activation(reg_activation_5_10), .reg_weight(reg_weight_5_10), .reg_partial_sum(reg_psum_5_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_11( .activation_in(reg_activation_5_10), .weight_in(reg_weight_4_11), .partial_sum_in(reg_psum_4_11), .reg_activation(reg_activation_5_11), .reg_weight(reg_weight_5_11), .reg_partial_sum(reg_psum_5_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_12( .activation_in(reg_activation_5_11), .weight_in(reg_weight_4_12), .partial_sum_in(reg_psum_4_12), .reg_activation(reg_activation_5_12), .reg_weight(reg_weight_5_12), .reg_partial_sum(reg_psum_5_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_13( .activation_in(reg_activation_5_12), .weight_in(reg_weight_4_13), .partial_sum_in(reg_psum_4_13), .reg_activation(reg_activation_5_13), .reg_weight(reg_weight_5_13), .reg_partial_sum(reg_psum_5_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_14( .activation_in(reg_activation_5_13), .weight_in(reg_weight_4_14), .partial_sum_in(reg_psum_4_14), .reg_activation(reg_activation_5_14), .reg_weight(reg_weight_5_14), .reg_partial_sum(reg_psum_5_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_15( .activation_in(reg_activation_5_14), .weight_in(reg_weight_4_15), .partial_sum_in(reg_psum_4_15), .reg_activation(reg_activation_5_15), .reg_weight(reg_weight_5_15), .reg_partial_sum(reg_psum_5_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_16( .activation_in(reg_activation_5_15), .weight_in(reg_weight_4_16), .partial_sum_in(reg_psum_4_16), .reg_activation(reg_activation_5_16), .reg_weight(reg_weight_5_16), .reg_partial_sum(reg_psum_5_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_17( .activation_in(reg_activation_5_16), .weight_in(reg_weight_4_17), .partial_sum_in(reg_psum_4_17), .reg_activation(reg_activation_5_17), .reg_weight(reg_weight_5_17), .reg_partial_sum(reg_psum_5_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_18( .activation_in(reg_activation_5_17), .weight_in(reg_weight_4_18), .partial_sum_in(reg_psum_4_18), .reg_activation(reg_activation_5_18), .reg_weight(reg_weight_5_18), .reg_partial_sum(reg_psum_5_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_19( .activation_in(reg_activation_5_18), .weight_in(reg_weight_4_19), .partial_sum_in(reg_psum_4_19), .reg_activation(reg_activation_5_19), .reg_weight(reg_weight_5_19), .reg_partial_sum(reg_psum_5_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_20( .activation_in(reg_activation_5_19), .weight_in(reg_weight_4_20), .partial_sum_in(reg_psum_4_20), .reg_activation(reg_activation_5_20), .reg_weight(reg_weight_5_20), .reg_partial_sum(reg_psum_5_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_21( .activation_in(reg_activation_5_20), .weight_in(reg_weight_4_21), .partial_sum_in(reg_psum_4_21), .reg_activation(reg_activation_5_21), .reg_weight(reg_weight_5_21), .reg_partial_sum(reg_psum_5_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_22( .activation_in(reg_activation_5_21), .weight_in(reg_weight_4_22), .partial_sum_in(reg_psum_4_22), .reg_activation(reg_activation_5_22), .reg_weight(reg_weight_5_22), .reg_partial_sum(reg_psum_5_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_23( .activation_in(reg_activation_5_22), .weight_in(reg_weight_4_23), .partial_sum_in(reg_psum_4_23), .reg_activation(reg_activation_5_23), .reg_weight(reg_weight_5_23), .reg_partial_sum(reg_psum_5_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_24( .activation_in(reg_activation_5_23), .weight_in(reg_weight_4_24), .partial_sum_in(reg_psum_4_24), .reg_activation(reg_activation_5_24), .reg_weight(reg_weight_5_24), .reg_partial_sum(reg_psum_5_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_25( .activation_in(reg_activation_5_24), .weight_in(reg_weight_4_25), .partial_sum_in(reg_psum_4_25), .reg_activation(reg_activation_5_25), .reg_weight(reg_weight_5_25), .reg_partial_sum(reg_psum_5_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_26( .activation_in(reg_activation_5_25), .weight_in(reg_weight_4_26), .partial_sum_in(reg_psum_4_26), .reg_activation(reg_activation_5_26), .reg_weight(reg_weight_5_26), .reg_partial_sum(reg_psum_5_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_27( .activation_in(reg_activation_5_26), .weight_in(reg_weight_4_27), .partial_sum_in(reg_psum_4_27), .reg_activation(reg_activation_5_27), .reg_weight(reg_weight_5_27), .reg_partial_sum(reg_psum_5_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_28( .activation_in(reg_activation_5_27), .weight_in(reg_weight_4_28), .partial_sum_in(reg_psum_4_28), .reg_activation(reg_activation_5_28), .reg_weight(reg_weight_5_28), .reg_partial_sum(reg_psum_5_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_29( .activation_in(reg_activation_5_28), .weight_in(reg_weight_4_29), .partial_sum_in(reg_psum_4_29), .reg_activation(reg_activation_5_29), .reg_weight(reg_weight_5_29), .reg_partial_sum(reg_psum_5_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_30( .activation_in(reg_activation_5_29), .weight_in(reg_weight_4_30), .partial_sum_in(reg_psum_4_30), .reg_activation(reg_activation_5_30), .reg_weight(reg_weight_5_30), .reg_partial_sum(reg_psum_5_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U5_31( .activation_in(reg_activation_5_30), .weight_in(reg_weight_4_31), .partial_sum_in(reg_psum_4_31), .reg_weight(reg_weight_5_31), .reg_partial_sum(reg_psum_5_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_0( .activation_in(in_activation_6), .weight_in(reg_weight_5_0), .partial_sum_in(reg_psum_5_0), .reg_activation(reg_activation_6_0), .reg_weight(reg_weight_6_0), .reg_partial_sum(reg_psum_6_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_1( .activation_in(reg_activation_6_0), .weight_in(reg_weight_5_1), .partial_sum_in(reg_psum_5_1), .reg_activation(reg_activation_6_1), .reg_weight(reg_weight_6_1), .reg_partial_sum(reg_psum_6_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_2( .activation_in(reg_activation_6_1), .weight_in(reg_weight_5_2), .partial_sum_in(reg_psum_5_2), .reg_activation(reg_activation_6_2), .reg_weight(reg_weight_6_2), .reg_partial_sum(reg_psum_6_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_3( .activation_in(reg_activation_6_2), .weight_in(reg_weight_5_3), .partial_sum_in(reg_psum_5_3), .reg_activation(reg_activation_6_3), .reg_weight(reg_weight_6_3), .reg_partial_sum(reg_psum_6_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_4( .activation_in(reg_activation_6_3), .weight_in(reg_weight_5_4), .partial_sum_in(reg_psum_5_4), .reg_activation(reg_activation_6_4), .reg_weight(reg_weight_6_4), .reg_partial_sum(reg_psum_6_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_5( .activation_in(reg_activation_6_4), .weight_in(reg_weight_5_5), .partial_sum_in(reg_psum_5_5), .reg_activation(reg_activation_6_5), .reg_weight(reg_weight_6_5), .reg_partial_sum(reg_psum_6_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_6( .activation_in(reg_activation_6_5), .weight_in(reg_weight_5_6), .partial_sum_in(reg_psum_5_6), .reg_activation(reg_activation_6_6), .reg_weight(reg_weight_6_6), .reg_partial_sum(reg_psum_6_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_7( .activation_in(reg_activation_6_6), .weight_in(reg_weight_5_7), .partial_sum_in(reg_psum_5_7), .reg_activation(reg_activation_6_7), .reg_weight(reg_weight_6_7), .reg_partial_sum(reg_psum_6_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_8( .activation_in(reg_activation_6_7), .weight_in(reg_weight_5_8), .partial_sum_in(reg_psum_5_8), .reg_activation(reg_activation_6_8), .reg_weight(reg_weight_6_8), .reg_partial_sum(reg_psum_6_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_9( .activation_in(reg_activation_6_8), .weight_in(reg_weight_5_9), .partial_sum_in(reg_psum_5_9), .reg_activation(reg_activation_6_9), .reg_weight(reg_weight_6_9), .reg_partial_sum(reg_psum_6_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_10( .activation_in(reg_activation_6_9), .weight_in(reg_weight_5_10), .partial_sum_in(reg_psum_5_10), .reg_activation(reg_activation_6_10), .reg_weight(reg_weight_6_10), .reg_partial_sum(reg_psum_6_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_11( .activation_in(reg_activation_6_10), .weight_in(reg_weight_5_11), .partial_sum_in(reg_psum_5_11), .reg_activation(reg_activation_6_11), .reg_weight(reg_weight_6_11), .reg_partial_sum(reg_psum_6_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_12( .activation_in(reg_activation_6_11), .weight_in(reg_weight_5_12), .partial_sum_in(reg_psum_5_12), .reg_activation(reg_activation_6_12), .reg_weight(reg_weight_6_12), .reg_partial_sum(reg_psum_6_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_13( .activation_in(reg_activation_6_12), .weight_in(reg_weight_5_13), .partial_sum_in(reg_psum_5_13), .reg_activation(reg_activation_6_13), .reg_weight(reg_weight_6_13), .reg_partial_sum(reg_psum_6_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_14( .activation_in(reg_activation_6_13), .weight_in(reg_weight_5_14), .partial_sum_in(reg_psum_5_14), .reg_activation(reg_activation_6_14), .reg_weight(reg_weight_6_14), .reg_partial_sum(reg_psum_6_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_15( .activation_in(reg_activation_6_14), .weight_in(reg_weight_5_15), .partial_sum_in(reg_psum_5_15), .reg_activation(reg_activation_6_15), .reg_weight(reg_weight_6_15), .reg_partial_sum(reg_psum_6_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_16( .activation_in(reg_activation_6_15), .weight_in(reg_weight_5_16), .partial_sum_in(reg_psum_5_16), .reg_activation(reg_activation_6_16), .reg_weight(reg_weight_6_16), .reg_partial_sum(reg_psum_6_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_17( .activation_in(reg_activation_6_16), .weight_in(reg_weight_5_17), .partial_sum_in(reg_psum_5_17), .reg_activation(reg_activation_6_17), .reg_weight(reg_weight_6_17), .reg_partial_sum(reg_psum_6_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_18( .activation_in(reg_activation_6_17), .weight_in(reg_weight_5_18), .partial_sum_in(reg_psum_5_18), .reg_activation(reg_activation_6_18), .reg_weight(reg_weight_6_18), .reg_partial_sum(reg_psum_6_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_19( .activation_in(reg_activation_6_18), .weight_in(reg_weight_5_19), .partial_sum_in(reg_psum_5_19), .reg_activation(reg_activation_6_19), .reg_weight(reg_weight_6_19), .reg_partial_sum(reg_psum_6_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_20( .activation_in(reg_activation_6_19), .weight_in(reg_weight_5_20), .partial_sum_in(reg_psum_5_20), .reg_activation(reg_activation_6_20), .reg_weight(reg_weight_6_20), .reg_partial_sum(reg_psum_6_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_21( .activation_in(reg_activation_6_20), .weight_in(reg_weight_5_21), .partial_sum_in(reg_psum_5_21), .reg_activation(reg_activation_6_21), .reg_weight(reg_weight_6_21), .reg_partial_sum(reg_psum_6_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_22( .activation_in(reg_activation_6_21), .weight_in(reg_weight_5_22), .partial_sum_in(reg_psum_5_22), .reg_activation(reg_activation_6_22), .reg_weight(reg_weight_6_22), .reg_partial_sum(reg_psum_6_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_23( .activation_in(reg_activation_6_22), .weight_in(reg_weight_5_23), .partial_sum_in(reg_psum_5_23), .reg_activation(reg_activation_6_23), .reg_weight(reg_weight_6_23), .reg_partial_sum(reg_psum_6_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_24( .activation_in(reg_activation_6_23), .weight_in(reg_weight_5_24), .partial_sum_in(reg_psum_5_24), .reg_activation(reg_activation_6_24), .reg_weight(reg_weight_6_24), .reg_partial_sum(reg_psum_6_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_25( .activation_in(reg_activation_6_24), .weight_in(reg_weight_5_25), .partial_sum_in(reg_psum_5_25), .reg_activation(reg_activation_6_25), .reg_weight(reg_weight_6_25), .reg_partial_sum(reg_psum_6_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_26( .activation_in(reg_activation_6_25), .weight_in(reg_weight_5_26), .partial_sum_in(reg_psum_5_26), .reg_activation(reg_activation_6_26), .reg_weight(reg_weight_6_26), .reg_partial_sum(reg_psum_6_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_27( .activation_in(reg_activation_6_26), .weight_in(reg_weight_5_27), .partial_sum_in(reg_psum_5_27), .reg_activation(reg_activation_6_27), .reg_weight(reg_weight_6_27), .reg_partial_sum(reg_psum_6_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_28( .activation_in(reg_activation_6_27), .weight_in(reg_weight_5_28), .partial_sum_in(reg_psum_5_28), .reg_activation(reg_activation_6_28), .reg_weight(reg_weight_6_28), .reg_partial_sum(reg_psum_6_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_29( .activation_in(reg_activation_6_28), .weight_in(reg_weight_5_29), .partial_sum_in(reg_psum_5_29), .reg_activation(reg_activation_6_29), .reg_weight(reg_weight_6_29), .reg_partial_sum(reg_psum_6_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_30( .activation_in(reg_activation_6_29), .weight_in(reg_weight_5_30), .partial_sum_in(fault_reg_psum_5_30), .reg_activation(reg_activation_6_30), .reg_weight(reg_weight_6_30), .reg_partial_sum(reg_psum_6_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U6_31( .activation_in(reg_activation_6_30), .weight_in(reg_weight_5_31), .partial_sum_in(reg_psum_5_31), .reg_weight(reg_weight_6_31), .reg_partial_sum(reg_psum_6_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_0( .activation_in(in_activation_7), .weight_in(reg_weight_6_0), .partial_sum_in(reg_psum_6_0), .reg_activation(reg_activation_7_0), .reg_weight(reg_weight_7_0), .reg_partial_sum(reg_psum_7_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_1( .activation_in(reg_activation_7_0), .weight_in(reg_weight_6_1), .partial_sum_in(reg_psum_6_1), .reg_activation(reg_activation_7_1), .reg_weight(reg_weight_7_1), .reg_partial_sum(reg_psum_7_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_2( .activation_in(reg_activation_7_1), .weight_in(reg_weight_6_2), .partial_sum_in(reg_psum_6_2), .reg_activation(reg_activation_7_2), .reg_weight(reg_weight_7_2), .reg_partial_sum(reg_psum_7_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_3( .activation_in(reg_activation_7_2), .weight_in(reg_weight_6_3), .partial_sum_in(reg_psum_6_3), .reg_activation(reg_activation_7_3), .reg_weight(reg_weight_7_3), .reg_partial_sum(reg_psum_7_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_4( .activation_in(reg_activation_7_3), .weight_in(reg_weight_6_4), .partial_sum_in(reg_psum_6_4), .reg_activation(reg_activation_7_4), .reg_weight(reg_weight_7_4), .reg_partial_sum(reg_psum_7_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_5( .activation_in(reg_activation_7_4), .weight_in(reg_weight_6_5), .partial_sum_in(reg_psum_6_5), .reg_activation(reg_activation_7_5), .reg_weight(reg_weight_7_5), .reg_partial_sum(reg_psum_7_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_6( .activation_in(reg_activation_7_5), .weight_in(reg_weight_6_6), .partial_sum_in(reg_psum_6_6), .reg_activation(reg_activation_7_6), .reg_weight(reg_weight_7_6), .reg_partial_sum(reg_psum_7_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_7( .activation_in(reg_activation_7_6), .weight_in(reg_weight_6_7), .partial_sum_in(reg_psum_6_7), .reg_activation(reg_activation_7_7), .reg_weight(reg_weight_7_7), .reg_partial_sum(reg_psum_7_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_8( .activation_in(reg_activation_7_7), .weight_in(reg_weight_6_8), .partial_sum_in(reg_psum_6_8), .reg_activation(reg_activation_7_8), .reg_weight(reg_weight_7_8), .reg_partial_sum(reg_psum_7_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_9( .activation_in(reg_activation_7_8), .weight_in(reg_weight_6_9), .partial_sum_in(reg_psum_6_9), .reg_activation(reg_activation_7_9), .reg_weight(reg_weight_7_9), .reg_partial_sum(reg_psum_7_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_10( .activation_in(reg_activation_7_9), .weight_in(reg_weight_6_10), .partial_sum_in(reg_psum_6_10), .reg_activation(reg_activation_7_10), .reg_weight(reg_weight_7_10), .reg_partial_sum(reg_psum_7_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_11( .activation_in(reg_activation_7_10), .weight_in(reg_weight_6_11), .partial_sum_in(reg_psum_6_11), .reg_activation(reg_activation_7_11), .reg_weight(reg_weight_7_11), .reg_partial_sum(reg_psum_7_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_12( .activation_in(reg_activation_7_11), .weight_in(reg_weight_6_12), .partial_sum_in(reg_psum_6_12), .reg_activation(reg_activation_7_12), .reg_weight(reg_weight_7_12), .reg_partial_sum(reg_psum_7_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_13( .activation_in(reg_activation_7_12), .weight_in(reg_weight_6_13), .partial_sum_in(reg_psum_6_13), .reg_activation(reg_activation_7_13), .reg_weight(reg_weight_7_13), .reg_partial_sum(reg_psum_7_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_14( .activation_in(reg_activation_7_13), .weight_in(reg_weight_6_14), .partial_sum_in(reg_psum_6_14), .reg_activation(reg_activation_7_14), .reg_weight(reg_weight_7_14), .reg_partial_sum(reg_psum_7_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_15( .activation_in(reg_activation_7_14), .weight_in(reg_weight_6_15), .partial_sum_in(reg_psum_6_15), .reg_activation(reg_activation_7_15), .reg_weight(reg_weight_7_15), .reg_partial_sum(reg_psum_7_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_16( .activation_in(reg_activation_7_15), .weight_in(reg_weight_6_16), .partial_sum_in(reg_psum_6_16), .reg_activation(reg_activation_7_16), .reg_weight(reg_weight_7_16), .reg_partial_sum(reg_psum_7_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_17( .activation_in(reg_activation_7_16), .weight_in(reg_weight_6_17), .partial_sum_in(reg_psum_6_17), .reg_activation(reg_activation_7_17), .reg_weight(reg_weight_7_17), .reg_partial_sum(reg_psum_7_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_18( .activation_in(reg_activation_7_17), .weight_in(reg_weight_6_18), .partial_sum_in(reg_psum_6_18), .reg_activation(reg_activation_7_18), .reg_weight(reg_weight_7_18), .reg_partial_sum(reg_psum_7_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_19( .activation_in(reg_activation_7_18), .weight_in(reg_weight_6_19), .partial_sum_in(reg_psum_6_19), .reg_activation(reg_activation_7_19), .reg_weight(reg_weight_7_19), .reg_partial_sum(reg_psum_7_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_20( .activation_in(reg_activation_7_19), .weight_in(reg_weight_6_20), .partial_sum_in(reg_psum_6_20), .reg_activation(reg_activation_7_20), .reg_weight(reg_weight_7_20), .reg_partial_sum(reg_psum_7_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_21( .activation_in(reg_activation_7_20), .weight_in(reg_weight_6_21), .partial_sum_in(reg_psum_6_21), .reg_activation(reg_activation_7_21), .reg_weight(reg_weight_7_21), .reg_partial_sum(reg_psum_7_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_22( .activation_in(reg_activation_7_21), .weight_in(reg_weight_6_22), .partial_sum_in(reg_psum_6_22), .reg_activation(reg_activation_7_22), .reg_weight(reg_weight_7_22), .reg_partial_sum(reg_psum_7_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_23( .activation_in(reg_activation_7_22), .weight_in(reg_weight_6_23), .partial_sum_in(reg_psum_6_23), .reg_activation(reg_activation_7_23), .reg_weight(reg_weight_7_23), .reg_partial_sum(reg_psum_7_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_24( .activation_in(reg_activation_7_23), .weight_in(reg_weight_6_24), .partial_sum_in(reg_psum_6_24), .reg_activation(reg_activation_7_24), .reg_weight(reg_weight_7_24), .reg_partial_sum(reg_psum_7_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_25( .activation_in(reg_activation_7_24), .weight_in(reg_weight_6_25), .partial_sum_in(reg_psum_6_25), .reg_activation(reg_activation_7_25), .reg_weight(reg_weight_7_25), .reg_partial_sum(reg_psum_7_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_26( .activation_in(reg_activation_7_25), .weight_in(reg_weight_6_26), .partial_sum_in(fault_reg_psum_6_26), .reg_activation(reg_activation_7_26), .reg_weight(reg_weight_7_26), .reg_partial_sum(reg_psum_7_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_27( .activation_in(reg_activation_7_26), .weight_in(reg_weight_6_27), .partial_sum_in(reg_psum_6_27), .reg_activation(reg_activation_7_27), .reg_weight(reg_weight_7_27), .reg_partial_sum(reg_psum_7_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_28( .activation_in(reg_activation_7_27), .weight_in(reg_weight_6_28), .partial_sum_in(reg_psum_6_28), .reg_activation(reg_activation_7_28), .reg_weight(reg_weight_7_28), .reg_partial_sum(reg_psum_7_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_29( .activation_in(reg_activation_7_28), .weight_in(reg_weight_6_29), .partial_sum_in(reg_psum_6_29), .reg_activation(reg_activation_7_29), .reg_weight(reg_weight_7_29), .reg_partial_sum(reg_psum_7_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_30( .activation_in(reg_activation_7_29), .weight_in(reg_weight_6_30), .partial_sum_in(reg_psum_6_30), .reg_activation(reg_activation_7_30), .reg_weight(reg_weight_7_30), .reg_partial_sum(reg_psum_7_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U7_31( .activation_in(reg_activation_7_30), .weight_in(reg_weight_6_31), .partial_sum_in(reg_psum_6_31), .reg_weight(reg_weight_7_31), .reg_partial_sum(reg_psum_7_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_0( .activation_in(in_activation_8), .weight_in(reg_weight_7_0), .partial_sum_in(reg_psum_7_0), .reg_activation(reg_activation_8_0), .reg_weight(reg_weight_8_0), .reg_partial_sum(reg_psum_8_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_1( .activation_in(reg_activation_8_0), .weight_in(reg_weight_7_1), .partial_sum_in(reg_psum_7_1), .reg_activation(reg_activation_8_1), .reg_weight(reg_weight_8_1), .reg_partial_sum(reg_psum_8_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_2( .activation_in(reg_activation_8_1), .weight_in(reg_weight_7_2), .partial_sum_in(reg_psum_7_2), .reg_activation(reg_activation_8_2), .reg_weight(reg_weight_8_2), .reg_partial_sum(reg_psum_8_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_3( .activation_in(reg_activation_8_2), .weight_in(reg_weight_7_3), .partial_sum_in(reg_psum_7_3), .reg_activation(reg_activation_8_3), .reg_weight(reg_weight_8_3), .reg_partial_sum(reg_psum_8_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_4( .activation_in(reg_activation_8_3), .weight_in(reg_weight_7_4), .partial_sum_in(reg_psum_7_4), .reg_activation(reg_activation_8_4), .reg_weight(reg_weight_8_4), .reg_partial_sum(reg_psum_8_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_5( .activation_in(reg_activation_8_4), .weight_in(reg_weight_7_5), .partial_sum_in(reg_psum_7_5), .reg_activation(reg_activation_8_5), .reg_weight(reg_weight_8_5), .reg_partial_sum(reg_psum_8_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_6( .activation_in(reg_activation_8_5), .weight_in(reg_weight_7_6), .partial_sum_in(reg_psum_7_6), .reg_activation(reg_activation_8_6), .reg_weight(reg_weight_8_6), .reg_partial_sum(reg_psum_8_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_7( .activation_in(reg_activation_8_6), .weight_in(reg_weight_7_7), .partial_sum_in(reg_psum_7_7), .reg_activation(reg_activation_8_7), .reg_weight(reg_weight_8_7), .reg_partial_sum(reg_psum_8_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_8( .activation_in(reg_activation_8_7), .weight_in(reg_weight_7_8), .partial_sum_in(reg_psum_7_8), .reg_activation(reg_activation_8_8), .reg_weight(reg_weight_8_8), .reg_partial_sum(reg_psum_8_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_9( .activation_in(reg_activation_8_8), .weight_in(reg_weight_7_9), .partial_sum_in(reg_psum_7_9), .reg_activation(reg_activation_8_9), .reg_weight(reg_weight_8_9), .reg_partial_sum(reg_psum_8_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_10( .activation_in(reg_activation_8_9), .weight_in(reg_weight_7_10), .partial_sum_in(reg_psum_7_10), .reg_activation(reg_activation_8_10), .reg_weight(reg_weight_8_10), .reg_partial_sum(reg_psum_8_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_11( .activation_in(reg_activation_8_10), .weight_in(reg_weight_7_11), .partial_sum_in(reg_psum_7_11), .reg_activation(reg_activation_8_11), .reg_weight(reg_weight_8_11), .reg_partial_sum(reg_psum_8_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_12( .activation_in(reg_activation_8_11), .weight_in(reg_weight_7_12), .partial_sum_in(reg_psum_7_12), .reg_activation(reg_activation_8_12), .reg_weight(reg_weight_8_12), .reg_partial_sum(reg_psum_8_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_13( .activation_in(reg_activation_8_12), .weight_in(reg_weight_7_13), .partial_sum_in(reg_psum_7_13), .reg_activation(reg_activation_8_13), .reg_weight(reg_weight_8_13), .reg_partial_sum(reg_psum_8_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_14( .activation_in(reg_activation_8_13), .weight_in(reg_weight_7_14), .partial_sum_in(reg_psum_7_14), .reg_activation(reg_activation_8_14), .reg_weight(reg_weight_8_14), .reg_partial_sum(reg_psum_8_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_15( .activation_in(reg_activation_8_14), .weight_in(reg_weight_7_15), .partial_sum_in(reg_psum_7_15), .reg_activation(reg_activation_8_15), .reg_weight(reg_weight_8_15), .reg_partial_sum(reg_psum_8_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_16( .activation_in(reg_activation_8_15), .weight_in(reg_weight_7_16), .partial_sum_in(reg_psum_7_16), .reg_activation(reg_activation_8_16), .reg_weight(reg_weight_8_16), .reg_partial_sum(reg_psum_8_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_17( .activation_in(reg_activation_8_16), .weight_in(reg_weight_7_17), .partial_sum_in(reg_psum_7_17), .reg_activation(reg_activation_8_17), .reg_weight(reg_weight_8_17), .reg_partial_sum(reg_psum_8_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_18( .activation_in(reg_activation_8_17), .weight_in(reg_weight_7_18), .partial_sum_in(reg_psum_7_18), .reg_activation(reg_activation_8_18), .reg_weight(reg_weight_8_18), .reg_partial_sum(reg_psum_8_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_19( .activation_in(reg_activation_8_18), .weight_in(reg_weight_7_19), .partial_sum_in(reg_psum_7_19), .reg_activation(reg_activation_8_19), .reg_weight(reg_weight_8_19), .reg_partial_sum(reg_psum_8_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_20( .activation_in(reg_activation_8_19), .weight_in(reg_weight_7_20), .partial_sum_in(reg_psum_7_20), .reg_activation(reg_activation_8_20), .reg_weight(reg_weight_8_20), .reg_partial_sum(reg_psum_8_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_21( .activation_in(reg_activation_8_20), .weight_in(reg_weight_7_21), .partial_sum_in(reg_psum_7_21), .reg_activation(reg_activation_8_21), .reg_weight(reg_weight_8_21), .reg_partial_sum(reg_psum_8_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_22( .activation_in(reg_activation_8_21), .weight_in(reg_weight_7_22), .partial_sum_in(reg_psum_7_22), .reg_activation(reg_activation_8_22), .reg_weight(reg_weight_8_22), .reg_partial_sum(reg_psum_8_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_23( .activation_in(reg_activation_8_22), .weight_in(reg_weight_7_23), .partial_sum_in(reg_psum_7_23), .reg_activation(reg_activation_8_23), .reg_weight(reg_weight_8_23), .reg_partial_sum(reg_psum_8_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_24( .activation_in(reg_activation_8_23), .weight_in(reg_weight_7_24), .partial_sum_in(reg_psum_7_24), .reg_activation(reg_activation_8_24), .reg_weight(reg_weight_8_24), .reg_partial_sum(reg_psum_8_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_25( .activation_in(reg_activation_8_24), .weight_in(reg_weight_7_25), .partial_sum_in(reg_psum_7_25), .reg_activation(reg_activation_8_25), .reg_weight(reg_weight_8_25), .reg_partial_sum(reg_psum_8_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_26( .activation_in(reg_activation_8_25), .weight_in(reg_weight_7_26), .partial_sum_in(reg_psum_7_26), .reg_activation(reg_activation_8_26), .reg_weight(reg_weight_8_26), .reg_partial_sum(reg_psum_8_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_27( .activation_in(reg_activation_8_26), .weight_in(reg_weight_7_27), .partial_sum_in(reg_psum_7_27), .reg_activation(reg_activation_8_27), .reg_weight(reg_weight_8_27), .reg_partial_sum(reg_psum_8_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_28( .activation_in(reg_activation_8_27), .weight_in(reg_weight_7_28), .partial_sum_in(reg_psum_7_28), .reg_activation(reg_activation_8_28), .reg_weight(reg_weight_8_28), .reg_partial_sum(reg_psum_8_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_29( .activation_in(reg_activation_8_28), .weight_in(reg_weight_7_29), .partial_sum_in(reg_psum_7_29), .reg_activation(reg_activation_8_29), .reg_weight(reg_weight_8_29), .reg_partial_sum(reg_psum_8_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_30( .activation_in(reg_activation_8_29), .weight_in(reg_weight_7_30), .partial_sum_in(reg_psum_7_30), .reg_activation(reg_activation_8_30), .reg_weight(reg_weight_8_30), .reg_partial_sum(reg_psum_8_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U8_31( .activation_in(reg_activation_8_30), .weight_in(reg_weight_7_31), .partial_sum_in(reg_psum_7_31), .reg_weight(reg_weight_8_31), .reg_partial_sum(reg_psum_8_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_0( .activation_in(in_activation_9), .weight_in(reg_weight_8_0), .partial_sum_in(reg_psum_8_0), .reg_activation(reg_activation_9_0), .reg_weight(reg_weight_9_0), .reg_partial_sum(reg_psum_9_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_1( .activation_in(reg_activation_9_0), .weight_in(reg_weight_8_1), .partial_sum_in(reg_psum_8_1), .reg_activation(reg_activation_9_1), .reg_weight(reg_weight_9_1), .reg_partial_sum(reg_psum_9_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_2( .activation_in(reg_activation_9_1), .weight_in(reg_weight_8_2), .partial_sum_in(reg_psum_8_2), .reg_activation(reg_activation_9_2), .reg_weight(reg_weight_9_2), .reg_partial_sum(reg_psum_9_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_3( .activation_in(reg_activation_9_2), .weight_in(reg_weight_8_3), .partial_sum_in(reg_psum_8_3), .reg_activation(reg_activation_9_3), .reg_weight(reg_weight_9_3), .reg_partial_sum(reg_psum_9_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_4( .activation_in(reg_activation_9_3), .weight_in(reg_weight_8_4), .partial_sum_in(reg_psum_8_4), .reg_activation(reg_activation_9_4), .reg_weight(reg_weight_9_4), .reg_partial_sum(reg_psum_9_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_5( .activation_in(reg_activation_9_4), .weight_in(reg_weight_8_5), .partial_sum_in(reg_psum_8_5), .reg_activation(reg_activation_9_5), .reg_weight(reg_weight_9_5), .reg_partial_sum(reg_psum_9_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_6( .activation_in(reg_activation_9_5), .weight_in(reg_weight_8_6), .partial_sum_in(reg_psum_8_6), .reg_activation(reg_activation_9_6), .reg_weight(reg_weight_9_6), .reg_partial_sum(reg_psum_9_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_7( .activation_in(reg_activation_9_6), .weight_in(reg_weight_8_7), .partial_sum_in(reg_psum_8_7), .reg_activation(reg_activation_9_7), .reg_weight(reg_weight_9_7), .reg_partial_sum(reg_psum_9_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_8( .activation_in(reg_activation_9_7), .weight_in(reg_weight_8_8), .partial_sum_in(reg_psum_8_8), .reg_activation(reg_activation_9_8), .reg_weight(reg_weight_9_8), .reg_partial_sum(reg_psum_9_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_9( .activation_in(reg_activation_9_8), .weight_in(reg_weight_8_9), .partial_sum_in(reg_psum_8_9), .reg_activation(reg_activation_9_9), .reg_weight(reg_weight_9_9), .reg_partial_sum(reg_psum_9_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_10( .activation_in(reg_activation_9_9), .weight_in(reg_weight_8_10), .partial_sum_in(reg_psum_8_10), .reg_activation(reg_activation_9_10), .reg_weight(reg_weight_9_10), .reg_partial_sum(reg_psum_9_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_11( .activation_in(reg_activation_9_10), .weight_in(reg_weight_8_11), .partial_sum_in(reg_psum_8_11), .reg_activation(reg_activation_9_11), .reg_weight(reg_weight_9_11), .reg_partial_sum(reg_psum_9_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_12( .activation_in(reg_activation_9_11), .weight_in(reg_weight_8_12), .partial_sum_in(reg_psum_8_12), .reg_activation(reg_activation_9_12), .reg_weight(reg_weight_9_12), .reg_partial_sum(reg_psum_9_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_13( .activation_in(reg_activation_9_12), .weight_in(reg_weight_8_13), .partial_sum_in(reg_psum_8_13), .reg_activation(reg_activation_9_13), .reg_weight(reg_weight_9_13), .reg_partial_sum(reg_psum_9_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_14( .activation_in(reg_activation_9_13), .weight_in(reg_weight_8_14), .partial_sum_in(reg_psum_8_14), .reg_activation(reg_activation_9_14), .reg_weight(reg_weight_9_14), .reg_partial_sum(reg_psum_9_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_15( .activation_in(reg_activation_9_14), .weight_in(reg_weight_8_15), .partial_sum_in(reg_psum_8_15), .reg_activation(reg_activation_9_15), .reg_weight(reg_weight_9_15), .reg_partial_sum(reg_psum_9_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_16( .activation_in(reg_activation_9_15), .weight_in(reg_weight_8_16), .partial_sum_in(reg_psum_8_16), .reg_activation(reg_activation_9_16), .reg_weight(reg_weight_9_16), .reg_partial_sum(reg_psum_9_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_17( .activation_in(reg_activation_9_16), .weight_in(reg_weight_8_17), .partial_sum_in(reg_psum_8_17), .reg_activation(reg_activation_9_17), .reg_weight(reg_weight_9_17), .reg_partial_sum(reg_psum_9_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_18( .activation_in(reg_activation_9_17), .weight_in(reg_weight_8_18), .partial_sum_in(reg_psum_8_18), .reg_activation(reg_activation_9_18), .reg_weight(reg_weight_9_18), .reg_partial_sum(reg_psum_9_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_19( .activation_in(reg_activation_9_18), .weight_in(reg_weight_8_19), .partial_sum_in(reg_psum_8_19), .reg_activation(reg_activation_9_19), .reg_weight(reg_weight_9_19), .reg_partial_sum(reg_psum_9_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_20( .activation_in(reg_activation_9_19), .weight_in(reg_weight_8_20), .partial_sum_in(reg_psum_8_20), .reg_activation(reg_activation_9_20), .reg_weight(reg_weight_9_20), .reg_partial_sum(reg_psum_9_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_21( .activation_in(reg_activation_9_20), .weight_in(reg_weight_8_21), .partial_sum_in(reg_psum_8_21), .reg_activation(reg_activation_9_21), .reg_weight(reg_weight_9_21), .reg_partial_sum(reg_psum_9_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_22( .activation_in(reg_activation_9_21), .weight_in(reg_weight_8_22), .partial_sum_in(reg_psum_8_22), .reg_activation(reg_activation_9_22), .reg_weight(reg_weight_9_22), .reg_partial_sum(reg_psum_9_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_23( .activation_in(reg_activation_9_22), .weight_in(reg_weight_8_23), .partial_sum_in(reg_psum_8_23), .reg_activation(reg_activation_9_23), .reg_weight(reg_weight_9_23), .reg_partial_sum(reg_psum_9_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_24( .activation_in(reg_activation_9_23), .weight_in(reg_weight_8_24), .partial_sum_in(reg_psum_8_24), .reg_activation(reg_activation_9_24), .reg_weight(reg_weight_9_24), .reg_partial_sum(reg_psum_9_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_25( .activation_in(reg_activation_9_24), .weight_in(reg_weight_8_25), .partial_sum_in(reg_psum_8_25), .reg_activation(reg_activation_9_25), .reg_weight(reg_weight_9_25), .reg_partial_sum(reg_psum_9_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_26( .activation_in(reg_activation_9_25), .weight_in(reg_weight_8_26), .partial_sum_in(reg_psum_8_26), .reg_activation(reg_activation_9_26), .reg_weight(reg_weight_9_26), .reg_partial_sum(reg_psum_9_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_27( .activation_in(reg_activation_9_26), .weight_in(reg_weight_8_27), .partial_sum_in(reg_psum_8_27), .reg_activation(reg_activation_9_27), .reg_weight(reg_weight_9_27), .reg_partial_sum(reg_psum_9_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_28( .activation_in(reg_activation_9_27), .weight_in(reg_weight_8_28), .partial_sum_in(reg_psum_8_28), .reg_activation(reg_activation_9_28), .reg_weight(reg_weight_9_28), .reg_partial_sum(reg_psum_9_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_29( .activation_in(reg_activation_9_28), .weight_in(reg_weight_8_29), .partial_sum_in(reg_psum_8_29), .reg_activation(reg_activation_9_29), .reg_weight(reg_weight_9_29), .reg_partial_sum(reg_psum_9_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_30( .activation_in(reg_activation_9_29), .weight_in(reg_weight_8_30), .partial_sum_in(reg_psum_8_30), .reg_activation(reg_activation_9_30), .reg_weight(reg_weight_9_30), .reg_partial_sum(reg_psum_9_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U9_31( .activation_in(reg_activation_9_30), .weight_in(reg_weight_8_31), .partial_sum_in(reg_psum_8_31), .reg_weight(reg_weight_9_31), .reg_partial_sum(reg_psum_9_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_0( .activation_in(in_activation_10), .weight_in(reg_weight_9_0), .partial_sum_in(reg_psum_9_0), .reg_activation(reg_activation_10_0), .reg_weight(reg_weight_10_0), .reg_partial_sum(reg_psum_10_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_1( .activation_in(reg_activation_10_0), .weight_in(reg_weight_9_1), .partial_sum_in(reg_psum_9_1), .reg_activation(reg_activation_10_1), .reg_weight(reg_weight_10_1), .reg_partial_sum(reg_psum_10_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_2( .activation_in(reg_activation_10_1), .weight_in(reg_weight_9_2), .partial_sum_in(reg_psum_9_2), .reg_activation(reg_activation_10_2), .reg_weight(reg_weight_10_2), .reg_partial_sum(reg_psum_10_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_3( .activation_in(reg_activation_10_2), .weight_in(reg_weight_9_3), .partial_sum_in(reg_psum_9_3), .reg_activation(reg_activation_10_3), .reg_weight(reg_weight_10_3), .reg_partial_sum(reg_psum_10_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_4( .activation_in(reg_activation_10_3), .weight_in(reg_weight_9_4), .partial_sum_in(reg_psum_9_4), .reg_activation(reg_activation_10_4), .reg_weight(reg_weight_10_4), .reg_partial_sum(reg_psum_10_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_5( .activation_in(reg_activation_10_4), .weight_in(reg_weight_9_5), .partial_sum_in(reg_psum_9_5), .reg_activation(reg_activation_10_5), .reg_weight(reg_weight_10_5), .reg_partial_sum(reg_psum_10_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_6( .activation_in(reg_activation_10_5), .weight_in(reg_weight_9_6), .partial_sum_in(reg_psum_9_6), .reg_activation(reg_activation_10_6), .reg_weight(reg_weight_10_6), .reg_partial_sum(reg_psum_10_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_7( .activation_in(reg_activation_10_6), .weight_in(reg_weight_9_7), .partial_sum_in(reg_psum_9_7), .reg_activation(reg_activation_10_7), .reg_weight(reg_weight_10_7), .reg_partial_sum(reg_psum_10_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_8( .activation_in(reg_activation_10_7), .weight_in(reg_weight_9_8), .partial_sum_in(reg_psum_9_8), .reg_activation(reg_activation_10_8), .reg_weight(reg_weight_10_8), .reg_partial_sum(reg_psum_10_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_9( .activation_in(reg_activation_10_8), .weight_in(reg_weight_9_9), .partial_sum_in(reg_psum_9_9), .reg_activation(reg_activation_10_9), .reg_weight(reg_weight_10_9), .reg_partial_sum(reg_psum_10_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_10( .activation_in(reg_activation_10_9), .weight_in(reg_weight_9_10), .partial_sum_in(reg_psum_9_10), .reg_activation(reg_activation_10_10), .reg_weight(reg_weight_10_10), .reg_partial_sum(reg_psum_10_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_11( .activation_in(reg_activation_10_10), .weight_in(reg_weight_9_11), .partial_sum_in(reg_psum_9_11), .reg_activation(reg_activation_10_11), .reg_weight(reg_weight_10_11), .reg_partial_sum(reg_psum_10_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_12( .activation_in(reg_activation_10_11), .weight_in(reg_weight_9_12), .partial_sum_in(reg_psum_9_12), .reg_activation(reg_activation_10_12), .reg_weight(reg_weight_10_12), .reg_partial_sum(reg_psum_10_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_13( .activation_in(reg_activation_10_12), .weight_in(reg_weight_9_13), .partial_sum_in(reg_psum_9_13), .reg_activation(reg_activation_10_13), .reg_weight(reg_weight_10_13), .reg_partial_sum(reg_psum_10_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_14( .activation_in(reg_activation_10_13), .weight_in(reg_weight_9_14), .partial_sum_in(reg_psum_9_14), .reg_activation(reg_activation_10_14), .reg_weight(reg_weight_10_14), .reg_partial_sum(reg_psum_10_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_15( .activation_in(reg_activation_10_14), .weight_in(reg_weight_9_15), .partial_sum_in(reg_psum_9_15), .reg_activation(reg_activation_10_15), .reg_weight(reg_weight_10_15), .reg_partial_sum(reg_psum_10_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_16( .activation_in(reg_activation_10_15), .weight_in(reg_weight_9_16), .partial_sum_in(reg_psum_9_16), .reg_activation(reg_activation_10_16), .reg_weight(reg_weight_10_16), .reg_partial_sum(reg_psum_10_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_17( .activation_in(reg_activation_10_16), .weight_in(reg_weight_9_17), .partial_sum_in(reg_psum_9_17), .reg_activation(reg_activation_10_17), .reg_weight(reg_weight_10_17), .reg_partial_sum(reg_psum_10_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_18( .activation_in(reg_activation_10_17), .weight_in(reg_weight_9_18), .partial_sum_in(reg_psum_9_18), .reg_activation(reg_activation_10_18), .reg_weight(reg_weight_10_18), .reg_partial_sum(reg_psum_10_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_19( .activation_in(reg_activation_10_18), .weight_in(reg_weight_9_19), .partial_sum_in(reg_psum_9_19), .reg_activation(reg_activation_10_19), .reg_weight(reg_weight_10_19), .reg_partial_sum(reg_psum_10_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_20( .activation_in(reg_activation_10_19), .weight_in(reg_weight_9_20), .partial_sum_in(reg_psum_9_20), .reg_activation(reg_activation_10_20), .reg_weight(reg_weight_10_20), .reg_partial_sum(reg_psum_10_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_21( .activation_in(reg_activation_10_20), .weight_in(reg_weight_9_21), .partial_sum_in(reg_psum_9_21), .reg_activation(reg_activation_10_21), .reg_weight(reg_weight_10_21), .reg_partial_sum(reg_psum_10_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_22( .activation_in(reg_activation_10_21), .weight_in(reg_weight_9_22), .partial_sum_in(reg_psum_9_22), .reg_activation(reg_activation_10_22), .reg_weight(reg_weight_10_22), .reg_partial_sum(reg_psum_10_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_23( .activation_in(reg_activation_10_22), .weight_in(reg_weight_9_23), .partial_sum_in(reg_psum_9_23), .reg_activation(reg_activation_10_23), .reg_weight(reg_weight_10_23), .reg_partial_sum(reg_psum_10_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_24( .activation_in(reg_activation_10_23), .weight_in(reg_weight_9_24), .partial_sum_in(reg_psum_9_24), .reg_activation(reg_activation_10_24), .reg_weight(reg_weight_10_24), .reg_partial_sum(reg_psum_10_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_25( .activation_in(reg_activation_10_24), .weight_in(reg_weight_9_25), .partial_sum_in(reg_psum_9_25), .reg_activation(reg_activation_10_25), .reg_weight(reg_weight_10_25), .reg_partial_sum(reg_psum_10_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_26( .activation_in(reg_activation_10_25), .weight_in(reg_weight_9_26), .partial_sum_in(reg_psum_9_26), .reg_activation(reg_activation_10_26), .reg_weight(reg_weight_10_26), .reg_partial_sum(reg_psum_10_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_27( .activation_in(reg_activation_10_26), .weight_in(reg_weight_9_27), .partial_sum_in(reg_psum_9_27), .reg_activation(reg_activation_10_27), .reg_weight(reg_weight_10_27), .reg_partial_sum(reg_psum_10_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_28( .activation_in(reg_activation_10_27), .weight_in(reg_weight_9_28), .partial_sum_in(reg_psum_9_28), .reg_activation(reg_activation_10_28), .reg_weight(reg_weight_10_28), .reg_partial_sum(reg_psum_10_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_29( .activation_in(reg_activation_10_28), .weight_in(reg_weight_9_29), .partial_sum_in(reg_psum_9_29), .reg_activation(reg_activation_10_29), .reg_weight(reg_weight_10_29), .reg_partial_sum(reg_psum_10_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_30( .activation_in(reg_activation_10_29), .weight_in(reg_weight_9_30), .partial_sum_in(reg_psum_9_30), .reg_activation(reg_activation_10_30), .reg_weight(reg_weight_10_30), .reg_partial_sum(reg_psum_10_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U10_31( .activation_in(reg_activation_10_30), .weight_in(reg_weight_9_31), .partial_sum_in(reg_psum_9_31), .reg_weight(reg_weight_10_31), .reg_partial_sum(reg_psum_10_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_0( .activation_in(in_activation_11), .weight_in(reg_weight_10_0), .partial_sum_in(reg_psum_10_0), .reg_activation(reg_activation_11_0), .reg_weight(reg_weight_11_0), .reg_partial_sum(reg_psum_11_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_1( .activation_in(reg_activation_11_0), .weight_in(reg_weight_10_1), .partial_sum_in(reg_psum_10_1), .reg_activation(reg_activation_11_1), .reg_weight(reg_weight_11_1), .reg_partial_sum(reg_psum_11_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_2( .activation_in(reg_activation_11_1), .weight_in(reg_weight_10_2), .partial_sum_in(reg_psum_10_2), .reg_activation(reg_activation_11_2), .reg_weight(reg_weight_11_2), .reg_partial_sum(reg_psum_11_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_3( .activation_in(reg_activation_11_2), .weight_in(reg_weight_10_3), .partial_sum_in(reg_psum_10_3), .reg_activation(reg_activation_11_3), .reg_weight(reg_weight_11_3), .reg_partial_sum(reg_psum_11_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_4( .activation_in(reg_activation_11_3), .weight_in(reg_weight_10_4), .partial_sum_in(reg_psum_10_4), .reg_activation(reg_activation_11_4), .reg_weight(reg_weight_11_4), .reg_partial_sum(reg_psum_11_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_5( .activation_in(reg_activation_11_4), .weight_in(reg_weight_10_5), .partial_sum_in(reg_psum_10_5), .reg_activation(reg_activation_11_5), .reg_weight(reg_weight_11_5), .reg_partial_sum(reg_psum_11_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_6( .activation_in(reg_activation_11_5), .weight_in(reg_weight_10_6), .partial_sum_in(reg_psum_10_6), .reg_activation(reg_activation_11_6), .reg_weight(reg_weight_11_6), .reg_partial_sum(reg_psum_11_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_7( .activation_in(reg_activation_11_6), .weight_in(reg_weight_10_7), .partial_sum_in(reg_psum_10_7), .reg_activation(reg_activation_11_7), .reg_weight(reg_weight_11_7), .reg_partial_sum(reg_psum_11_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_8( .activation_in(reg_activation_11_7), .weight_in(reg_weight_10_8), .partial_sum_in(reg_psum_10_8), .reg_activation(reg_activation_11_8), .reg_weight(reg_weight_11_8), .reg_partial_sum(reg_psum_11_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_9( .activation_in(reg_activation_11_8), .weight_in(reg_weight_10_9), .partial_sum_in(reg_psum_10_9), .reg_activation(reg_activation_11_9), .reg_weight(reg_weight_11_9), .reg_partial_sum(reg_psum_11_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_10( .activation_in(reg_activation_11_9), .weight_in(reg_weight_10_10), .partial_sum_in(reg_psum_10_10), .reg_activation(reg_activation_11_10), .reg_weight(reg_weight_11_10), .reg_partial_sum(reg_psum_11_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_11( .activation_in(reg_activation_11_10), .weight_in(reg_weight_10_11), .partial_sum_in(reg_psum_10_11), .reg_activation(reg_activation_11_11), .reg_weight(reg_weight_11_11), .reg_partial_sum(reg_psum_11_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_12( .activation_in(reg_activation_11_11), .weight_in(reg_weight_10_12), .partial_sum_in(reg_psum_10_12), .reg_activation(reg_activation_11_12), .reg_weight(reg_weight_11_12), .reg_partial_sum(reg_psum_11_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_13( .activation_in(reg_activation_11_12), .weight_in(reg_weight_10_13), .partial_sum_in(reg_psum_10_13), .reg_activation(reg_activation_11_13), .reg_weight(reg_weight_11_13), .reg_partial_sum(reg_psum_11_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_14( .activation_in(reg_activation_11_13), .weight_in(reg_weight_10_14), .partial_sum_in(reg_psum_10_14), .reg_activation(reg_activation_11_14), .reg_weight(reg_weight_11_14), .reg_partial_sum(reg_psum_11_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_15( .activation_in(reg_activation_11_14), .weight_in(reg_weight_10_15), .partial_sum_in(reg_psum_10_15), .reg_activation(reg_activation_11_15), .reg_weight(reg_weight_11_15), .reg_partial_sum(reg_psum_11_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_16( .activation_in(reg_activation_11_15), .weight_in(reg_weight_10_16), .partial_sum_in(reg_psum_10_16), .reg_activation(reg_activation_11_16), .reg_weight(reg_weight_11_16), .reg_partial_sum(reg_psum_11_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_17( .activation_in(reg_activation_11_16), .weight_in(reg_weight_10_17), .partial_sum_in(reg_psum_10_17), .reg_activation(reg_activation_11_17), .reg_weight(reg_weight_11_17), .reg_partial_sum(reg_psum_11_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_18( .activation_in(reg_activation_11_17), .weight_in(reg_weight_10_18), .partial_sum_in(reg_psum_10_18), .reg_activation(reg_activation_11_18), .reg_weight(reg_weight_11_18), .reg_partial_sum(reg_psum_11_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_19( .activation_in(reg_activation_11_18), .weight_in(reg_weight_10_19), .partial_sum_in(reg_psum_10_19), .reg_activation(reg_activation_11_19), .reg_weight(reg_weight_11_19), .reg_partial_sum(reg_psum_11_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_20( .activation_in(reg_activation_11_19), .weight_in(reg_weight_10_20), .partial_sum_in(reg_psum_10_20), .reg_activation(reg_activation_11_20), .reg_weight(reg_weight_11_20), .reg_partial_sum(reg_psum_11_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_21( .activation_in(reg_activation_11_20), .weight_in(reg_weight_10_21), .partial_sum_in(reg_psum_10_21), .reg_activation(reg_activation_11_21), .reg_weight(reg_weight_11_21), .reg_partial_sum(reg_psum_11_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_22( .activation_in(reg_activation_11_21), .weight_in(reg_weight_10_22), .partial_sum_in(reg_psum_10_22), .reg_activation(reg_activation_11_22), .reg_weight(reg_weight_11_22), .reg_partial_sum(reg_psum_11_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_23( .activation_in(reg_activation_11_22), .weight_in(reg_weight_10_23), .partial_sum_in(reg_psum_10_23), .reg_activation(reg_activation_11_23), .reg_weight(reg_weight_11_23), .reg_partial_sum(reg_psum_11_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_24( .activation_in(reg_activation_11_23), .weight_in(reg_weight_10_24), .partial_sum_in(reg_psum_10_24), .reg_activation(reg_activation_11_24), .reg_weight(reg_weight_11_24), .reg_partial_sum(reg_psum_11_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_25( .activation_in(reg_activation_11_24), .weight_in(reg_weight_10_25), .partial_sum_in(reg_psum_10_25), .reg_activation(reg_activation_11_25), .reg_weight(reg_weight_11_25), .reg_partial_sum(reg_psum_11_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_26( .activation_in(reg_activation_11_25), .weight_in(reg_weight_10_26), .partial_sum_in(fault_reg_psum_10_26), .reg_activation(reg_activation_11_26), .reg_weight(reg_weight_11_26), .reg_partial_sum(reg_psum_11_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_27( .activation_in(reg_activation_11_26), .weight_in(reg_weight_10_27), .partial_sum_in(reg_psum_10_27), .reg_activation(reg_activation_11_27), .reg_weight(reg_weight_11_27), .reg_partial_sum(reg_psum_11_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_28( .activation_in(reg_activation_11_27), .weight_in(reg_weight_10_28), .partial_sum_in(reg_psum_10_28), .reg_activation(reg_activation_11_28), .reg_weight(reg_weight_11_28), .reg_partial_sum(reg_psum_11_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_29( .activation_in(reg_activation_11_28), .weight_in(reg_weight_10_29), .partial_sum_in(reg_psum_10_29), .reg_activation(reg_activation_11_29), .reg_weight(reg_weight_11_29), .reg_partial_sum(reg_psum_11_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_30( .activation_in(reg_activation_11_29), .weight_in(reg_weight_10_30), .partial_sum_in(reg_psum_10_30), .reg_activation(reg_activation_11_30), .reg_weight(reg_weight_11_30), .reg_partial_sum(reg_psum_11_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U11_31( .activation_in(reg_activation_11_30), .weight_in(reg_weight_10_31), .partial_sum_in(reg_psum_10_31), .reg_weight(reg_weight_11_31), .reg_partial_sum(reg_psum_11_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_0( .activation_in(in_activation_12), .weight_in(reg_weight_11_0), .partial_sum_in(reg_psum_11_0), .reg_activation(reg_activation_12_0), .reg_weight(reg_weight_12_0), .reg_partial_sum(reg_psum_12_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_1( .activation_in(reg_activation_12_0), .weight_in(reg_weight_11_1), .partial_sum_in(reg_psum_11_1), .reg_activation(reg_activation_12_1), .reg_weight(reg_weight_12_1), .reg_partial_sum(reg_psum_12_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_2( .activation_in(reg_activation_12_1), .weight_in(reg_weight_11_2), .partial_sum_in(reg_psum_11_2), .reg_activation(reg_activation_12_2), .reg_weight(reg_weight_12_2), .reg_partial_sum(reg_psum_12_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_3( .activation_in(reg_activation_12_2), .weight_in(reg_weight_11_3), .partial_sum_in(reg_psum_11_3), .reg_activation(reg_activation_12_3), .reg_weight(reg_weight_12_3), .reg_partial_sum(reg_psum_12_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_4( .activation_in(reg_activation_12_3), .weight_in(reg_weight_11_4), .partial_sum_in(reg_psum_11_4), .reg_activation(reg_activation_12_4), .reg_weight(reg_weight_12_4), .reg_partial_sum(reg_psum_12_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_5( .activation_in(reg_activation_12_4), .weight_in(reg_weight_11_5), .partial_sum_in(reg_psum_11_5), .reg_activation(reg_activation_12_5), .reg_weight(reg_weight_12_5), .reg_partial_sum(reg_psum_12_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_6( .activation_in(reg_activation_12_5), .weight_in(reg_weight_11_6), .partial_sum_in(reg_psum_11_6), .reg_activation(reg_activation_12_6), .reg_weight(reg_weight_12_6), .reg_partial_sum(reg_psum_12_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_7( .activation_in(reg_activation_12_6), .weight_in(reg_weight_11_7), .partial_sum_in(reg_psum_11_7), .reg_activation(reg_activation_12_7), .reg_weight(reg_weight_12_7), .reg_partial_sum(reg_psum_12_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_8( .activation_in(reg_activation_12_7), .weight_in(reg_weight_11_8), .partial_sum_in(reg_psum_11_8), .reg_activation(reg_activation_12_8), .reg_weight(reg_weight_12_8), .reg_partial_sum(reg_psum_12_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_9( .activation_in(reg_activation_12_8), .weight_in(reg_weight_11_9), .partial_sum_in(reg_psum_11_9), .reg_activation(reg_activation_12_9), .reg_weight(reg_weight_12_9), .reg_partial_sum(reg_psum_12_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_10( .activation_in(reg_activation_12_9), .weight_in(reg_weight_11_10), .partial_sum_in(reg_psum_11_10), .reg_activation(reg_activation_12_10), .reg_weight(reg_weight_12_10), .reg_partial_sum(reg_psum_12_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_11( .activation_in(reg_activation_12_10), .weight_in(reg_weight_11_11), .partial_sum_in(reg_psum_11_11), .reg_activation(reg_activation_12_11), .reg_weight(reg_weight_12_11), .reg_partial_sum(reg_psum_12_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_12( .activation_in(reg_activation_12_11), .weight_in(reg_weight_11_12), .partial_sum_in(reg_psum_11_12), .reg_activation(reg_activation_12_12), .reg_weight(reg_weight_12_12), .reg_partial_sum(reg_psum_12_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_13( .activation_in(reg_activation_12_12), .weight_in(reg_weight_11_13), .partial_sum_in(reg_psum_11_13), .reg_activation(reg_activation_12_13), .reg_weight(reg_weight_12_13), .reg_partial_sum(reg_psum_12_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_14( .activation_in(reg_activation_12_13), .weight_in(reg_weight_11_14), .partial_sum_in(reg_psum_11_14), .reg_activation(reg_activation_12_14), .reg_weight(reg_weight_12_14), .reg_partial_sum(reg_psum_12_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_15( .activation_in(reg_activation_12_14), .weight_in(reg_weight_11_15), .partial_sum_in(reg_psum_11_15), .reg_activation(reg_activation_12_15), .reg_weight(reg_weight_12_15), .reg_partial_sum(reg_psum_12_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_16( .activation_in(reg_activation_12_15), .weight_in(reg_weight_11_16), .partial_sum_in(reg_psum_11_16), .reg_activation(reg_activation_12_16), .reg_weight(reg_weight_12_16), .reg_partial_sum(reg_psum_12_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_17( .activation_in(reg_activation_12_16), .weight_in(reg_weight_11_17), .partial_sum_in(reg_psum_11_17), .reg_activation(reg_activation_12_17), .reg_weight(reg_weight_12_17), .reg_partial_sum(reg_psum_12_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_18( .activation_in(reg_activation_12_17), .weight_in(reg_weight_11_18), .partial_sum_in(reg_psum_11_18), .reg_activation(reg_activation_12_18), .reg_weight(reg_weight_12_18), .reg_partial_sum(reg_psum_12_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_19( .activation_in(reg_activation_12_18), .weight_in(reg_weight_11_19), .partial_sum_in(reg_psum_11_19), .reg_activation(reg_activation_12_19), .reg_weight(reg_weight_12_19), .reg_partial_sum(reg_psum_12_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_20( .activation_in(reg_activation_12_19), .weight_in(reg_weight_11_20), .partial_sum_in(reg_psum_11_20), .reg_activation(reg_activation_12_20), .reg_weight(reg_weight_12_20), .reg_partial_sum(reg_psum_12_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_21( .activation_in(reg_activation_12_20), .weight_in(reg_weight_11_21), .partial_sum_in(reg_psum_11_21), .reg_activation(reg_activation_12_21), .reg_weight(reg_weight_12_21), .reg_partial_sum(reg_psum_12_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_22( .activation_in(reg_activation_12_21), .weight_in(reg_weight_11_22), .partial_sum_in(reg_psum_11_22), .reg_activation(reg_activation_12_22), .reg_weight(reg_weight_12_22), .reg_partial_sum(reg_psum_12_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_23( .activation_in(reg_activation_12_22), .weight_in(reg_weight_11_23), .partial_sum_in(reg_psum_11_23), .reg_activation(reg_activation_12_23), .reg_weight(reg_weight_12_23), .reg_partial_sum(reg_psum_12_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_24( .activation_in(reg_activation_12_23), .weight_in(reg_weight_11_24), .partial_sum_in(reg_psum_11_24), .reg_activation(reg_activation_12_24), .reg_weight(reg_weight_12_24), .reg_partial_sum(reg_psum_12_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_25( .activation_in(reg_activation_12_24), .weight_in(reg_weight_11_25), .partial_sum_in(reg_psum_11_25), .reg_activation(reg_activation_12_25), .reg_weight(reg_weight_12_25), .reg_partial_sum(reg_psum_12_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_26( .activation_in(reg_activation_12_25), .weight_in(reg_weight_11_26), .partial_sum_in(reg_psum_11_26), .reg_activation(reg_activation_12_26), .reg_weight(reg_weight_12_26), .reg_partial_sum(reg_psum_12_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_27( .activation_in(reg_activation_12_26), .weight_in(reg_weight_11_27), .partial_sum_in(reg_psum_11_27), .reg_activation(reg_activation_12_27), .reg_weight(reg_weight_12_27), .reg_partial_sum(reg_psum_12_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_28( .activation_in(reg_activation_12_27), .weight_in(reg_weight_11_28), .partial_sum_in(reg_psum_11_28), .reg_activation(reg_activation_12_28), .reg_weight(reg_weight_12_28), .reg_partial_sum(reg_psum_12_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_29( .activation_in(reg_activation_12_28), .weight_in(reg_weight_11_29), .partial_sum_in(reg_psum_11_29), .reg_activation(reg_activation_12_29), .reg_weight(reg_weight_12_29), .reg_partial_sum(reg_psum_12_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_30( .activation_in(reg_activation_12_29), .weight_in(reg_weight_11_30), .partial_sum_in(reg_psum_11_30), .reg_activation(reg_activation_12_30), .reg_weight(reg_weight_12_30), .reg_partial_sum(reg_psum_12_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U12_31( .activation_in(reg_activation_12_30), .weight_in(reg_weight_11_31), .partial_sum_in(reg_psum_11_31), .reg_weight(reg_weight_12_31), .reg_partial_sum(reg_psum_12_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_0( .activation_in(in_activation_13), .weight_in(reg_weight_12_0), .partial_sum_in(reg_psum_12_0), .reg_activation(reg_activation_13_0), .reg_weight(reg_weight_13_0), .reg_partial_sum(reg_psum_13_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_1( .activation_in(reg_activation_13_0), .weight_in(reg_weight_12_1), .partial_sum_in(reg_psum_12_1), .reg_activation(reg_activation_13_1), .reg_weight(reg_weight_13_1), .reg_partial_sum(reg_psum_13_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_2( .activation_in(reg_activation_13_1), .weight_in(reg_weight_12_2), .partial_sum_in(reg_psum_12_2), .reg_activation(reg_activation_13_2), .reg_weight(reg_weight_13_2), .reg_partial_sum(reg_psum_13_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_3( .activation_in(reg_activation_13_2), .weight_in(reg_weight_12_3), .partial_sum_in(reg_psum_12_3), .reg_activation(reg_activation_13_3), .reg_weight(reg_weight_13_3), .reg_partial_sum(reg_psum_13_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_4( .activation_in(reg_activation_13_3), .weight_in(reg_weight_12_4), .partial_sum_in(reg_psum_12_4), .reg_activation(reg_activation_13_4), .reg_weight(reg_weight_13_4), .reg_partial_sum(reg_psum_13_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_5( .activation_in(reg_activation_13_4), .weight_in(reg_weight_12_5), .partial_sum_in(reg_psum_12_5), .reg_activation(reg_activation_13_5), .reg_weight(reg_weight_13_5), .reg_partial_sum(reg_psum_13_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_6( .activation_in(reg_activation_13_5), .weight_in(reg_weight_12_6), .partial_sum_in(reg_psum_12_6), .reg_activation(reg_activation_13_6), .reg_weight(reg_weight_13_6), .reg_partial_sum(reg_psum_13_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_7( .activation_in(reg_activation_13_6), .weight_in(reg_weight_12_7), .partial_sum_in(reg_psum_12_7), .reg_activation(reg_activation_13_7), .reg_weight(reg_weight_13_7), .reg_partial_sum(reg_psum_13_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_8( .activation_in(reg_activation_13_7), .weight_in(reg_weight_12_8), .partial_sum_in(reg_psum_12_8), .reg_activation(reg_activation_13_8), .reg_weight(reg_weight_13_8), .reg_partial_sum(reg_psum_13_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_9( .activation_in(reg_activation_13_8), .weight_in(reg_weight_12_9), .partial_sum_in(reg_psum_12_9), .reg_activation(reg_activation_13_9), .reg_weight(reg_weight_13_9), .reg_partial_sum(reg_psum_13_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_10( .activation_in(reg_activation_13_9), .weight_in(reg_weight_12_10), .partial_sum_in(reg_psum_12_10), .reg_activation(reg_activation_13_10), .reg_weight(reg_weight_13_10), .reg_partial_sum(reg_psum_13_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_11( .activation_in(reg_activation_13_10), .weight_in(reg_weight_12_11), .partial_sum_in(reg_psum_12_11), .reg_activation(reg_activation_13_11), .reg_weight(reg_weight_13_11), .reg_partial_sum(reg_psum_13_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_12( .activation_in(reg_activation_13_11), .weight_in(reg_weight_12_12), .partial_sum_in(reg_psum_12_12), .reg_activation(reg_activation_13_12), .reg_weight(reg_weight_13_12), .reg_partial_sum(reg_psum_13_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_13( .activation_in(reg_activation_13_12), .weight_in(reg_weight_12_13), .partial_sum_in(reg_psum_12_13), .reg_activation(reg_activation_13_13), .reg_weight(reg_weight_13_13), .reg_partial_sum(reg_psum_13_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_14( .activation_in(reg_activation_13_13), .weight_in(reg_weight_12_14), .partial_sum_in(reg_psum_12_14), .reg_activation(reg_activation_13_14), .reg_weight(reg_weight_13_14), .reg_partial_sum(reg_psum_13_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_15( .activation_in(reg_activation_13_14), .weight_in(reg_weight_12_15), .partial_sum_in(reg_psum_12_15), .reg_activation(reg_activation_13_15), .reg_weight(reg_weight_13_15), .reg_partial_sum(reg_psum_13_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_16( .activation_in(reg_activation_13_15), .weight_in(reg_weight_12_16), .partial_sum_in(reg_psum_12_16), .reg_activation(reg_activation_13_16), .reg_weight(reg_weight_13_16), .reg_partial_sum(reg_psum_13_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_17( .activation_in(reg_activation_13_16), .weight_in(reg_weight_12_17), .partial_sum_in(reg_psum_12_17), .reg_activation(reg_activation_13_17), .reg_weight(reg_weight_13_17), .reg_partial_sum(reg_psum_13_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_18( .activation_in(reg_activation_13_17), .weight_in(reg_weight_12_18), .partial_sum_in(reg_psum_12_18), .reg_activation(reg_activation_13_18), .reg_weight(reg_weight_13_18), .reg_partial_sum(reg_psum_13_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_19( .activation_in(reg_activation_13_18), .weight_in(reg_weight_12_19), .partial_sum_in(reg_psum_12_19), .reg_activation(reg_activation_13_19), .reg_weight(reg_weight_13_19), .reg_partial_sum(reg_psum_13_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_20( .activation_in(reg_activation_13_19), .weight_in(reg_weight_12_20), .partial_sum_in(reg_psum_12_20), .reg_activation(reg_activation_13_20), .reg_weight(reg_weight_13_20), .reg_partial_sum(reg_psum_13_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_21( .activation_in(reg_activation_13_20), .weight_in(reg_weight_12_21), .partial_sum_in(reg_psum_12_21), .reg_activation(reg_activation_13_21), .reg_weight(reg_weight_13_21), .reg_partial_sum(reg_psum_13_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_22( .activation_in(reg_activation_13_21), .weight_in(reg_weight_12_22), .partial_sum_in(reg_psum_12_22), .reg_activation(reg_activation_13_22), .reg_weight(reg_weight_13_22), .reg_partial_sum(reg_psum_13_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_23( .activation_in(reg_activation_13_22), .weight_in(reg_weight_12_23), .partial_sum_in(reg_psum_12_23), .reg_activation(reg_activation_13_23), .reg_weight(reg_weight_13_23), .reg_partial_sum(reg_psum_13_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_24( .activation_in(reg_activation_13_23), .weight_in(reg_weight_12_24), .partial_sum_in(reg_psum_12_24), .reg_activation(reg_activation_13_24), .reg_weight(reg_weight_13_24), .reg_partial_sum(reg_psum_13_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_25( .activation_in(reg_activation_13_24), .weight_in(reg_weight_12_25), .partial_sum_in(reg_psum_12_25), .reg_activation(reg_activation_13_25), .reg_weight(reg_weight_13_25), .reg_partial_sum(reg_psum_13_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_26( .activation_in(reg_activation_13_25), .weight_in(reg_weight_12_26), .partial_sum_in(reg_psum_12_26), .reg_activation(reg_activation_13_26), .reg_weight(reg_weight_13_26), .reg_partial_sum(reg_psum_13_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_27( .activation_in(reg_activation_13_26), .weight_in(reg_weight_12_27), .partial_sum_in(reg_psum_12_27), .reg_activation(reg_activation_13_27), .reg_weight(reg_weight_13_27), .reg_partial_sum(reg_psum_13_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_28( .activation_in(reg_activation_13_27), .weight_in(reg_weight_12_28), .partial_sum_in(reg_psum_12_28), .reg_activation(reg_activation_13_28), .reg_weight(reg_weight_13_28), .reg_partial_sum(reg_psum_13_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_29( .activation_in(reg_activation_13_28), .weight_in(reg_weight_12_29), .partial_sum_in(reg_psum_12_29), .reg_activation(reg_activation_13_29), .reg_weight(reg_weight_13_29), .reg_partial_sum(reg_psum_13_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_30( .activation_in(reg_activation_13_29), .weight_in(reg_weight_12_30), .partial_sum_in(reg_psum_12_30), .reg_activation(reg_activation_13_30), .reg_weight(reg_weight_13_30), .reg_partial_sum(reg_psum_13_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U13_31( .activation_in(reg_activation_13_30), .weight_in(reg_weight_12_31), .partial_sum_in(reg_psum_12_31), .reg_weight(reg_weight_13_31), .reg_partial_sum(reg_psum_13_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_0( .activation_in(in_activation_14), .weight_in(reg_weight_13_0), .partial_sum_in(reg_psum_13_0), .reg_activation(reg_activation_14_0), .reg_weight(reg_weight_14_0), .reg_partial_sum(reg_psum_14_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_1( .activation_in(reg_activation_14_0), .weight_in(reg_weight_13_1), .partial_sum_in(reg_psum_13_1), .reg_activation(reg_activation_14_1), .reg_weight(reg_weight_14_1), .reg_partial_sum(reg_psum_14_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_2( .activation_in(reg_activation_14_1), .weight_in(reg_weight_13_2), .partial_sum_in(reg_psum_13_2), .reg_activation(reg_activation_14_2), .reg_weight(reg_weight_14_2), .reg_partial_sum(reg_psum_14_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_3( .activation_in(reg_activation_14_2), .weight_in(reg_weight_13_3), .partial_sum_in(fault_reg_psum_13_3), .reg_activation(reg_activation_14_3), .reg_weight(reg_weight_14_3), .reg_partial_sum(reg_psum_14_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_4( .activation_in(reg_activation_14_3), .weight_in(reg_weight_13_4), .partial_sum_in(reg_psum_13_4), .reg_activation(reg_activation_14_4), .reg_weight(reg_weight_14_4), .reg_partial_sum(reg_psum_14_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_5( .activation_in(reg_activation_14_4), .weight_in(reg_weight_13_5), .partial_sum_in(reg_psum_13_5), .reg_activation(reg_activation_14_5), .reg_weight(reg_weight_14_5), .reg_partial_sum(reg_psum_14_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_6( .activation_in(reg_activation_14_5), .weight_in(reg_weight_13_6), .partial_sum_in(reg_psum_13_6), .reg_activation(reg_activation_14_6), .reg_weight(reg_weight_14_6), .reg_partial_sum(reg_psum_14_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_7( .activation_in(reg_activation_14_6), .weight_in(reg_weight_13_7), .partial_sum_in(reg_psum_13_7), .reg_activation(reg_activation_14_7), .reg_weight(reg_weight_14_7), .reg_partial_sum(reg_psum_14_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_8( .activation_in(reg_activation_14_7), .weight_in(reg_weight_13_8), .partial_sum_in(reg_psum_13_8), .reg_activation(reg_activation_14_8), .reg_weight(reg_weight_14_8), .reg_partial_sum(reg_psum_14_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_9( .activation_in(reg_activation_14_8), .weight_in(reg_weight_13_9), .partial_sum_in(reg_psum_13_9), .reg_activation(reg_activation_14_9), .reg_weight(reg_weight_14_9), .reg_partial_sum(reg_psum_14_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_10( .activation_in(reg_activation_14_9), .weight_in(reg_weight_13_10), .partial_sum_in(reg_psum_13_10), .reg_activation(reg_activation_14_10), .reg_weight(reg_weight_14_10), .reg_partial_sum(reg_psum_14_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_11( .activation_in(reg_activation_14_10), .weight_in(reg_weight_13_11), .partial_sum_in(reg_psum_13_11), .reg_activation(reg_activation_14_11), .reg_weight(reg_weight_14_11), .reg_partial_sum(reg_psum_14_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_12( .activation_in(reg_activation_14_11), .weight_in(reg_weight_13_12), .partial_sum_in(reg_psum_13_12), .reg_activation(reg_activation_14_12), .reg_weight(reg_weight_14_12), .reg_partial_sum(reg_psum_14_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_13( .activation_in(reg_activation_14_12), .weight_in(reg_weight_13_13), .partial_sum_in(reg_psum_13_13), .reg_activation(reg_activation_14_13), .reg_weight(reg_weight_14_13), .reg_partial_sum(reg_psum_14_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_14( .activation_in(reg_activation_14_13), .weight_in(reg_weight_13_14), .partial_sum_in(reg_psum_13_14), .reg_activation(reg_activation_14_14), .reg_weight(reg_weight_14_14), .reg_partial_sum(reg_psum_14_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_15( .activation_in(reg_activation_14_14), .weight_in(reg_weight_13_15), .partial_sum_in(reg_psum_13_15), .reg_activation(reg_activation_14_15), .reg_weight(reg_weight_14_15), .reg_partial_sum(reg_psum_14_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_16( .activation_in(reg_activation_14_15), .weight_in(reg_weight_13_16), .partial_sum_in(reg_psum_13_16), .reg_activation(reg_activation_14_16), .reg_weight(reg_weight_14_16), .reg_partial_sum(reg_psum_14_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_17( .activation_in(reg_activation_14_16), .weight_in(reg_weight_13_17), .partial_sum_in(reg_psum_13_17), .reg_activation(reg_activation_14_17), .reg_weight(reg_weight_14_17), .reg_partial_sum(reg_psum_14_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_18( .activation_in(reg_activation_14_17), .weight_in(reg_weight_13_18), .partial_sum_in(reg_psum_13_18), .reg_activation(reg_activation_14_18), .reg_weight(reg_weight_14_18), .reg_partial_sum(reg_psum_14_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_19( .activation_in(reg_activation_14_18), .weight_in(reg_weight_13_19), .partial_sum_in(reg_psum_13_19), .reg_activation(reg_activation_14_19), .reg_weight(reg_weight_14_19), .reg_partial_sum(reg_psum_14_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_20( .activation_in(reg_activation_14_19), .weight_in(reg_weight_13_20), .partial_sum_in(reg_psum_13_20), .reg_activation(reg_activation_14_20), .reg_weight(reg_weight_14_20), .reg_partial_sum(reg_psum_14_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_21( .activation_in(reg_activation_14_20), .weight_in(reg_weight_13_21), .partial_sum_in(reg_psum_13_21), .reg_activation(reg_activation_14_21), .reg_weight(reg_weight_14_21), .reg_partial_sum(reg_psum_14_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_22( .activation_in(reg_activation_14_21), .weight_in(reg_weight_13_22), .partial_sum_in(reg_psum_13_22), .reg_activation(reg_activation_14_22), .reg_weight(reg_weight_14_22), .reg_partial_sum(reg_psum_14_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_23( .activation_in(reg_activation_14_22), .weight_in(reg_weight_13_23), .partial_sum_in(reg_psum_13_23), .reg_activation(reg_activation_14_23), .reg_weight(reg_weight_14_23), .reg_partial_sum(reg_psum_14_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_24( .activation_in(reg_activation_14_23), .weight_in(reg_weight_13_24), .partial_sum_in(reg_psum_13_24), .reg_activation(reg_activation_14_24), .reg_weight(reg_weight_14_24), .reg_partial_sum(reg_psum_14_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_25( .activation_in(reg_activation_14_24), .weight_in(reg_weight_13_25), .partial_sum_in(reg_psum_13_25), .reg_activation(reg_activation_14_25), .reg_weight(reg_weight_14_25), .reg_partial_sum(reg_psum_14_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_26( .activation_in(reg_activation_14_25), .weight_in(reg_weight_13_26), .partial_sum_in(reg_psum_13_26), .reg_activation(reg_activation_14_26), .reg_weight(reg_weight_14_26), .reg_partial_sum(reg_psum_14_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_27( .activation_in(reg_activation_14_26), .weight_in(reg_weight_13_27), .partial_sum_in(reg_psum_13_27), .reg_activation(reg_activation_14_27), .reg_weight(reg_weight_14_27), .reg_partial_sum(reg_psum_14_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_28( .activation_in(reg_activation_14_27), .weight_in(reg_weight_13_28), .partial_sum_in(reg_psum_13_28), .reg_activation(reg_activation_14_28), .reg_weight(reg_weight_14_28), .reg_partial_sum(reg_psum_14_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_29( .activation_in(reg_activation_14_28), .weight_in(reg_weight_13_29), .partial_sum_in(reg_psum_13_29), .reg_activation(reg_activation_14_29), .reg_weight(reg_weight_14_29), .reg_partial_sum(reg_psum_14_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_30( .activation_in(reg_activation_14_29), .weight_in(reg_weight_13_30), .partial_sum_in(reg_psum_13_30), .reg_activation(reg_activation_14_30), .reg_weight(reg_weight_14_30), .reg_partial_sum(reg_psum_14_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U14_31( .activation_in(reg_activation_14_30), .weight_in(reg_weight_13_31), .partial_sum_in(reg_psum_13_31), .reg_weight(reg_weight_14_31), .reg_partial_sum(reg_psum_14_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_0( .activation_in(in_activation_15), .weight_in(reg_weight_14_0), .partial_sum_in(reg_psum_14_0), .reg_activation(reg_activation_15_0), .reg_weight(reg_weight_15_0), .reg_partial_sum(reg_psum_15_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_1( .activation_in(reg_activation_15_0), .weight_in(reg_weight_14_1), .partial_sum_in(reg_psum_14_1), .reg_activation(reg_activation_15_1), .reg_weight(reg_weight_15_1), .reg_partial_sum(reg_psum_15_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_2( .activation_in(reg_activation_15_1), .weight_in(reg_weight_14_2), .partial_sum_in(reg_psum_14_2), .reg_activation(reg_activation_15_2), .reg_weight(reg_weight_15_2), .reg_partial_sum(reg_psum_15_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_3( .activation_in(reg_activation_15_2), .weight_in(reg_weight_14_3), .partial_sum_in(reg_psum_14_3), .reg_activation(reg_activation_15_3), .reg_weight(reg_weight_15_3), .reg_partial_sum(reg_psum_15_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_4( .activation_in(reg_activation_15_3), .weight_in(reg_weight_14_4), .partial_sum_in(reg_psum_14_4), .reg_activation(reg_activation_15_4), .reg_weight(reg_weight_15_4), .reg_partial_sum(reg_psum_15_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_5( .activation_in(reg_activation_15_4), .weight_in(reg_weight_14_5), .partial_sum_in(reg_psum_14_5), .reg_activation(reg_activation_15_5), .reg_weight(reg_weight_15_5), .reg_partial_sum(reg_psum_15_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_6( .activation_in(reg_activation_15_5), .weight_in(reg_weight_14_6), .partial_sum_in(reg_psum_14_6), .reg_activation(reg_activation_15_6), .reg_weight(reg_weight_15_6), .reg_partial_sum(reg_psum_15_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_7( .activation_in(reg_activation_15_6), .weight_in(reg_weight_14_7), .partial_sum_in(reg_psum_14_7), .reg_activation(reg_activation_15_7), .reg_weight(reg_weight_15_7), .reg_partial_sum(reg_psum_15_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_8( .activation_in(reg_activation_15_7), .weight_in(reg_weight_14_8), .partial_sum_in(reg_psum_14_8), .reg_activation(reg_activation_15_8), .reg_weight(reg_weight_15_8), .reg_partial_sum(reg_psum_15_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_9( .activation_in(reg_activation_15_8), .weight_in(reg_weight_14_9), .partial_sum_in(reg_psum_14_9), .reg_activation(reg_activation_15_9), .reg_weight(reg_weight_15_9), .reg_partial_sum(reg_psum_15_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_10( .activation_in(reg_activation_15_9), .weight_in(reg_weight_14_10), .partial_sum_in(reg_psum_14_10), .reg_activation(reg_activation_15_10), .reg_weight(reg_weight_15_10), .reg_partial_sum(reg_psum_15_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_11( .activation_in(reg_activation_15_10), .weight_in(reg_weight_14_11), .partial_sum_in(reg_psum_14_11), .reg_activation(reg_activation_15_11), .reg_weight(reg_weight_15_11), .reg_partial_sum(reg_psum_15_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_12( .activation_in(reg_activation_15_11), .weight_in(reg_weight_14_12), .partial_sum_in(reg_psum_14_12), .reg_activation(reg_activation_15_12), .reg_weight(reg_weight_15_12), .reg_partial_sum(reg_psum_15_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_13( .activation_in(reg_activation_15_12), .weight_in(reg_weight_14_13), .partial_sum_in(reg_psum_14_13), .reg_activation(reg_activation_15_13), .reg_weight(reg_weight_15_13), .reg_partial_sum(reg_psum_15_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_14( .activation_in(reg_activation_15_13), .weight_in(reg_weight_14_14), .partial_sum_in(reg_psum_14_14), .reg_activation(reg_activation_15_14), .reg_weight(reg_weight_15_14), .reg_partial_sum(reg_psum_15_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_15( .activation_in(reg_activation_15_14), .weight_in(reg_weight_14_15), .partial_sum_in(reg_psum_14_15), .reg_activation(reg_activation_15_15), .reg_weight(reg_weight_15_15), .reg_partial_sum(reg_psum_15_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_16( .activation_in(reg_activation_15_15), .weight_in(reg_weight_14_16), .partial_sum_in(reg_psum_14_16), .reg_activation(reg_activation_15_16), .reg_weight(reg_weight_15_16), .reg_partial_sum(reg_psum_15_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_17( .activation_in(reg_activation_15_16), .weight_in(reg_weight_14_17), .partial_sum_in(reg_psum_14_17), .reg_activation(reg_activation_15_17), .reg_weight(reg_weight_15_17), .reg_partial_sum(reg_psum_15_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_18( .activation_in(reg_activation_15_17), .weight_in(reg_weight_14_18), .partial_sum_in(reg_psum_14_18), .reg_activation(reg_activation_15_18), .reg_weight(reg_weight_15_18), .reg_partial_sum(reg_psum_15_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_19( .activation_in(reg_activation_15_18), .weight_in(reg_weight_14_19), .partial_sum_in(reg_psum_14_19), .reg_activation(reg_activation_15_19), .reg_weight(reg_weight_15_19), .reg_partial_sum(reg_psum_15_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_20( .activation_in(reg_activation_15_19), .weight_in(reg_weight_14_20), .partial_sum_in(fault_reg_psum_14_20), .reg_activation(reg_activation_15_20), .reg_weight(reg_weight_15_20), .reg_partial_sum(reg_psum_15_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_21( .activation_in(reg_activation_15_20), .weight_in(reg_weight_14_21), .partial_sum_in(reg_psum_14_21), .reg_activation(reg_activation_15_21), .reg_weight(reg_weight_15_21), .reg_partial_sum(reg_psum_15_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_22( .activation_in(reg_activation_15_21), .weight_in(reg_weight_14_22), .partial_sum_in(reg_psum_14_22), .reg_activation(reg_activation_15_22), .reg_weight(reg_weight_15_22), .reg_partial_sum(reg_psum_15_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_23( .activation_in(reg_activation_15_22), .weight_in(reg_weight_14_23), .partial_sum_in(reg_psum_14_23), .reg_activation(reg_activation_15_23), .reg_weight(reg_weight_15_23), .reg_partial_sum(reg_psum_15_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_24( .activation_in(reg_activation_15_23), .weight_in(reg_weight_14_24), .partial_sum_in(reg_psum_14_24), .reg_activation(reg_activation_15_24), .reg_weight(reg_weight_15_24), .reg_partial_sum(reg_psum_15_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_25( .activation_in(reg_activation_15_24), .weight_in(reg_weight_14_25), .partial_sum_in(reg_psum_14_25), .reg_activation(reg_activation_15_25), .reg_weight(reg_weight_15_25), .reg_partial_sum(reg_psum_15_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_26( .activation_in(reg_activation_15_25), .weight_in(reg_weight_14_26), .partial_sum_in(reg_psum_14_26), .reg_activation(reg_activation_15_26), .reg_weight(reg_weight_15_26), .reg_partial_sum(reg_psum_15_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_27( .activation_in(reg_activation_15_26), .weight_in(reg_weight_14_27), .partial_sum_in(reg_psum_14_27), .reg_activation(reg_activation_15_27), .reg_weight(reg_weight_15_27), .reg_partial_sum(reg_psum_15_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_28( .activation_in(reg_activation_15_27), .weight_in(reg_weight_14_28), .partial_sum_in(reg_psum_14_28), .reg_activation(reg_activation_15_28), .reg_weight(reg_weight_15_28), .reg_partial_sum(reg_psum_15_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_29( .activation_in(reg_activation_15_28), .weight_in(reg_weight_14_29), .partial_sum_in(reg_psum_14_29), .reg_activation(reg_activation_15_29), .reg_weight(reg_weight_15_29), .reg_partial_sum(reg_psum_15_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_30( .activation_in(reg_activation_15_29), .weight_in(reg_weight_14_30), .partial_sum_in(reg_psum_14_30), .reg_activation(reg_activation_15_30), .reg_weight(reg_weight_15_30), .reg_partial_sum(reg_psum_15_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U15_31( .activation_in(reg_activation_15_30), .weight_in(reg_weight_14_31), .partial_sum_in(reg_psum_14_31), .reg_weight(reg_weight_15_31), .reg_partial_sum(reg_psum_15_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_0( .activation_in(in_activation_16), .weight_in(reg_weight_15_0), .partial_sum_in(reg_psum_15_0), .reg_activation(reg_activation_16_0), .reg_weight(reg_weight_16_0), .reg_partial_sum(reg_psum_16_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_1( .activation_in(reg_activation_16_0), .weight_in(reg_weight_15_1), .partial_sum_in(reg_psum_15_1), .reg_activation(reg_activation_16_1), .reg_weight(reg_weight_16_1), .reg_partial_sum(reg_psum_16_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_2( .activation_in(reg_activation_16_1), .weight_in(reg_weight_15_2), .partial_sum_in(reg_psum_15_2), .reg_activation(reg_activation_16_2), .reg_weight(reg_weight_16_2), .reg_partial_sum(reg_psum_16_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_3( .activation_in(reg_activation_16_2), .weight_in(reg_weight_15_3), .partial_sum_in(reg_psum_15_3), .reg_activation(reg_activation_16_3), .reg_weight(reg_weight_16_3), .reg_partial_sum(reg_psum_16_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_4( .activation_in(reg_activation_16_3), .weight_in(reg_weight_15_4), .partial_sum_in(reg_psum_15_4), .reg_activation(reg_activation_16_4), .reg_weight(reg_weight_16_4), .reg_partial_sum(reg_psum_16_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_5( .activation_in(reg_activation_16_4), .weight_in(reg_weight_15_5), .partial_sum_in(reg_psum_15_5), .reg_activation(reg_activation_16_5), .reg_weight(reg_weight_16_5), .reg_partial_sum(reg_psum_16_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_6( .activation_in(reg_activation_16_5), .weight_in(reg_weight_15_6), .partial_sum_in(reg_psum_15_6), .reg_activation(reg_activation_16_6), .reg_weight(reg_weight_16_6), .reg_partial_sum(reg_psum_16_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_7( .activation_in(reg_activation_16_6), .weight_in(reg_weight_15_7), .partial_sum_in(reg_psum_15_7), .reg_activation(reg_activation_16_7), .reg_weight(reg_weight_16_7), .reg_partial_sum(reg_psum_16_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_8( .activation_in(reg_activation_16_7), .weight_in(reg_weight_15_8), .partial_sum_in(reg_psum_15_8), .reg_activation(reg_activation_16_8), .reg_weight(reg_weight_16_8), .reg_partial_sum(reg_psum_16_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_9( .activation_in(reg_activation_16_8), .weight_in(reg_weight_15_9), .partial_sum_in(reg_psum_15_9), .reg_activation(reg_activation_16_9), .reg_weight(reg_weight_16_9), .reg_partial_sum(reg_psum_16_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_10( .activation_in(reg_activation_16_9), .weight_in(reg_weight_15_10), .partial_sum_in(reg_psum_15_10), .reg_activation(reg_activation_16_10), .reg_weight(reg_weight_16_10), .reg_partial_sum(reg_psum_16_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_11( .activation_in(reg_activation_16_10), .weight_in(reg_weight_15_11), .partial_sum_in(reg_psum_15_11), .reg_activation(reg_activation_16_11), .reg_weight(reg_weight_16_11), .reg_partial_sum(reg_psum_16_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_12( .activation_in(reg_activation_16_11), .weight_in(reg_weight_15_12), .partial_sum_in(reg_psum_15_12), .reg_activation(reg_activation_16_12), .reg_weight(reg_weight_16_12), .reg_partial_sum(reg_psum_16_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_13( .activation_in(reg_activation_16_12), .weight_in(reg_weight_15_13), .partial_sum_in(reg_psum_15_13), .reg_activation(reg_activation_16_13), .reg_weight(reg_weight_16_13), .reg_partial_sum(reg_psum_16_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_14( .activation_in(reg_activation_16_13), .weight_in(reg_weight_15_14), .partial_sum_in(reg_psum_15_14), .reg_activation(reg_activation_16_14), .reg_weight(reg_weight_16_14), .reg_partial_sum(reg_psum_16_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_15( .activation_in(reg_activation_16_14), .weight_in(reg_weight_15_15), .partial_sum_in(reg_psum_15_15), .reg_activation(reg_activation_16_15), .reg_weight(reg_weight_16_15), .reg_partial_sum(reg_psum_16_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_16( .activation_in(reg_activation_16_15), .weight_in(reg_weight_15_16), .partial_sum_in(reg_psum_15_16), .reg_activation(reg_activation_16_16), .reg_weight(reg_weight_16_16), .reg_partial_sum(reg_psum_16_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_17( .activation_in(reg_activation_16_16), .weight_in(reg_weight_15_17), .partial_sum_in(reg_psum_15_17), .reg_activation(reg_activation_16_17), .reg_weight(reg_weight_16_17), .reg_partial_sum(reg_psum_16_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_18( .activation_in(reg_activation_16_17), .weight_in(reg_weight_15_18), .partial_sum_in(reg_psum_15_18), .reg_activation(reg_activation_16_18), .reg_weight(reg_weight_16_18), .reg_partial_sum(reg_psum_16_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_19( .activation_in(reg_activation_16_18), .weight_in(reg_weight_15_19), .partial_sum_in(reg_psum_15_19), .reg_activation(reg_activation_16_19), .reg_weight(reg_weight_16_19), .reg_partial_sum(reg_psum_16_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_20( .activation_in(reg_activation_16_19), .weight_in(reg_weight_15_20), .partial_sum_in(reg_psum_15_20), .reg_activation(reg_activation_16_20), .reg_weight(reg_weight_16_20), .reg_partial_sum(reg_psum_16_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_21( .activation_in(reg_activation_16_20), .weight_in(reg_weight_15_21), .partial_sum_in(reg_psum_15_21), .reg_activation(reg_activation_16_21), .reg_weight(reg_weight_16_21), .reg_partial_sum(reg_psum_16_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_22( .activation_in(reg_activation_16_21), .weight_in(reg_weight_15_22), .partial_sum_in(reg_psum_15_22), .reg_activation(reg_activation_16_22), .reg_weight(reg_weight_16_22), .reg_partial_sum(reg_psum_16_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_23( .activation_in(reg_activation_16_22), .weight_in(reg_weight_15_23), .partial_sum_in(reg_psum_15_23), .reg_activation(reg_activation_16_23), .reg_weight(reg_weight_16_23), .reg_partial_sum(reg_psum_16_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_24( .activation_in(reg_activation_16_23), .weight_in(reg_weight_15_24), .partial_sum_in(reg_psum_15_24), .reg_activation(reg_activation_16_24), .reg_weight(reg_weight_16_24), .reg_partial_sum(reg_psum_16_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_25( .activation_in(reg_activation_16_24), .weight_in(reg_weight_15_25), .partial_sum_in(reg_psum_15_25), .reg_activation(reg_activation_16_25), .reg_weight(reg_weight_16_25), .reg_partial_sum(reg_psum_16_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_26( .activation_in(reg_activation_16_25), .weight_in(reg_weight_15_26), .partial_sum_in(reg_psum_15_26), .reg_activation(reg_activation_16_26), .reg_weight(reg_weight_16_26), .reg_partial_sum(reg_psum_16_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_27( .activation_in(reg_activation_16_26), .weight_in(reg_weight_15_27), .partial_sum_in(reg_psum_15_27), .reg_activation(reg_activation_16_27), .reg_weight(reg_weight_16_27), .reg_partial_sum(reg_psum_16_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_28( .activation_in(reg_activation_16_27), .weight_in(reg_weight_15_28), .partial_sum_in(reg_psum_15_28), .reg_activation(reg_activation_16_28), .reg_weight(reg_weight_16_28), .reg_partial_sum(reg_psum_16_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_29( .activation_in(reg_activation_16_28), .weight_in(reg_weight_15_29), .partial_sum_in(reg_psum_15_29), .reg_activation(reg_activation_16_29), .reg_weight(reg_weight_16_29), .reg_partial_sum(reg_psum_16_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_30( .activation_in(reg_activation_16_29), .weight_in(reg_weight_15_30), .partial_sum_in(reg_psum_15_30), .reg_activation(reg_activation_16_30), .reg_weight(reg_weight_16_30), .reg_partial_sum(reg_psum_16_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U16_31( .activation_in(reg_activation_16_30), .weight_in(reg_weight_15_31), .partial_sum_in(reg_psum_15_31), .reg_weight(reg_weight_16_31), .reg_partial_sum(reg_psum_16_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_0( .activation_in(in_activation_17), .weight_in(reg_weight_16_0), .partial_sum_in(reg_psum_16_0), .reg_activation(reg_activation_17_0), .reg_weight(reg_weight_17_0), .reg_partial_sum(reg_psum_17_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_1( .activation_in(reg_activation_17_0), .weight_in(reg_weight_16_1), .partial_sum_in(reg_psum_16_1), .reg_activation(reg_activation_17_1), .reg_weight(reg_weight_17_1), .reg_partial_sum(reg_psum_17_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_2( .activation_in(reg_activation_17_1), .weight_in(reg_weight_16_2), .partial_sum_in(reg_psum_16_2), .reg_activation(reg_activation_17_2), .reg_weight(reg_weight_17_2), .reg_partial_sum(reg_psum_17_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_3( .activation_in(reg_activation_17_2), .weight_in(reg_weight_16_3), .partial_sum_in(reg_psum_16_3), .reg_activation(reg_activation_17_3), .reg_weight(reg_weight_17_3), .reg_partial_sum(reg_psum_17_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_4( .activation_in(reg_activation_17_3), .weight_in(reg_weight_16_4), .partial_sum_in(reg_psum_16_4), .reg_activation(reg_activation_17_4), .reg_weight(reg_weight_17_4), .reg_partial_sum(reg_psum_17_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_5( .activation_in(reg_activation_17_4), .weight_in(reg_weight_16_5), .partial_sum_in(fault_reg_psum_16_5), .reg_activation(reg_activation_17_5), .reg_weight(reg_weight_17_5), .reg_partial_sum(reg_psum_17_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_6( .activation_in(reg_activation_17_5), .weight_in(reg_weight_16_6), .partial_sum_in(reg_psum_16_6), .reg_activation(reg_activation_17_6), .reg_weight(reg_weight_17_6), .reg_partial_sum(reg_psum_17_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_7( .activation_in(reg_activation_17_6), .weight_in(reg_weight_16_7), .partial_sum_in(reg_psum_16_7), .reg_activation(reg_activation_17_7), .reg_weight(reg_weight_17_7), .reg_partial_sum(reg_psum_17_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_8( .activation_in(reg_activation_17_7), .weight_in(reg_weight_16_8), .partial_sum_in(reg_psum_16_8), .reg_activation(reg_activation_17_8), .reg_weight(reg_weight_17_8), .reg_partial_sum(reg_psum_17_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_9( .activation_in(reg_activation_17_8), .weight_in(reg_weight_16_9), .partial_sum_in(reg_psum_16_9), .reg_activation(reg_activation_17_9), .reg_weight(reg_weight_17_9), .reg_partial_sum(reg_psum_17_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_10( .activation_in(reg_activation_17_9), .weight_in(reg_weight_16_10), .partial_sum_in(reg_psum_16_10), .reg_activation(reg_activation_17_10), .reg_weight(reg_weight_17_10), .reg_partial_sum(reg_psum_17_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_11( .activation_in(reg_activation_17_10), .weight_in(reg_weight_16_11), .partial_sum_in(reg_psum_16_11), .reg_activation(reg_activation_17_11), .reg_weight(reg_weight_17_11), .reg_partial_sum(reg_psum_17_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_12( .activation_in(reg_activation_17_11), .weight_in(reg_weight_16_12), .partial_sum_in(reg_psum_16_12), .reg_activation(reg_activation_17_12), .reg_weight(reg_weight_17_12), .reg_partial_sum(reg_psum_17_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_13( .activation_in(reg_activation_17_12), .weight_in(reg_weight_16_13), .partial_sum_in(reg_psum_16_13), .reg_activation(reg_activation_17_13), .reg_weight(reg_weight_17_13), .reg_partial_sum(reg_psum_17_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_14( .activation_in(reg_activation_17_13), .weight_in(reg_weight_16_14), .partial_sum_in(reg_psum_16_14), .reg_activation(reg_activation_17_14), .reg_weight(reg_weight_17_14), .reg_partial_sum(reg_psum_17_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_15( .activation_in(reg_activation_17_14), .weight_in(reg_weight_16_15), .partial_sum_in(reg_psum_16_15), .reg_activation(reg_activation_17_15), .reg_weight(reg_weight_17_15), .reg_partial_sum(reg_psum_17_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_16( .activation_in(reg_activation_17_15), .weight_in(reg_weight_16_16), .partial_sum_in(reg_psum_16_16), .reg_activation(reg_activation_17_16), .reg_weight(reg_weight_17_16), .reg_partial_sum(reg_psum_17_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_17( .activation_in(reg_activation_17_16), .weight_in(reg_weight_16_17), .partial_sum_in(reg_psum_16_17), .reg_activation(reg_activation_17_17), .reg_weight(reg_weight_17_17), .reg_partial_sum(reg_psum_17_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_18( .activation_in(reg_activation_17_17), .weight_in(reg_weight_16_18), .partial_sum_in(reg_psum_16_18), .reg_activation(reg_activation_17_18), .reg_weight(reg_weight_17_18), .reg_partial_sum(reg_psum_17_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_19( .activation_in(reg_activation_17_18), .weight_in(reg_weight_16_19), .partial_sum_in(reg_psum_16_19), .reg_activation(reg_activation_17_19), .reg_weight(reg_weight_17_19), .reg_partial_sum(reg_psum_17_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_20( .activation_in(reg_activation_17_19), .weight_in(reg_weight_16_20), .partial_sum_in(reg_psum_16_20), .reg_activation(reg_activation_17_20), .reg_weight(reg_weight_17_20), .reg_partial_sum(reg_psum_17_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_21( .activation_in(reg_activation_17_20), .weight_in(reg_weight_16_21), .partial_sum_in(reg_psum_16_21), .reg_activation(reg_activation_17_21), .reg_weight(reg_weight_17_21), .reg_partial_sum(reg_psum_17_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_22( .activation_in(reg_activation_17_21), .weight_in(reg_weight_16_22), .partial_sum_in(reg_psum_16_22), .reg_activation(reg_activation_17_22), .reg_weight(reg_weight_17_22), .reg_partial_sum(reg_psum_17_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_23( .activation_in(reg_activation_17_22), .weight_in(reg_weight_16_23), .partial_sum_in(reg_psum_16_23), .reg_activation(reg_activation_17_23), .reg_weight(reg_weight_17_23), .reg_partial_sum(reg_psum_17_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_24( .activation_in(reg_activation_17_23), .weight_in(reg_weight_16_24), .partial_sum_in(reg_psum_16_24), .reg_activation(reg_activation_17_24), .reg_weight(reg_weight_17_24), .reg_partial_sum(reg_psum_17_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_25( .activation_in(reg_activation_17_24), .weight_in(reg_weight_16_25), .partial_sum_in(reg_psum_16_25), .reg_activation(reg_activation_17_25), .reg_weight(reg_weight_17_25), .reg_partial_sum(reg_psum_17_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_26( .activation_in(reg_activation_17_25), .weight_in(reg_weight_16_26), .partial_sum_in(reg_psum_16_26), .reg_activation(reg_activation_17_26), .reg_weight(reg_weight_17_26), .reg_partial_sum(reg_psum_17_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_27( .activation_in(reg_activation_17_26), .weight_in(reg_weight_16_27), .partial_sum_in(reg_psum_16_27), .reg_activation(reg_activation_17_27), .reg_weight(reg_weight_17_27), .reg_partial_sum(reg_psum_17_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_28( .activation_in(reg_activation_17_27), .weight_in(reg_weight_16_28), .partial_sum_in(reg_psum_16_28), .reg_activation(reg_activation_17_28), .reg_weight(reg_weight_17_28), .reg_partial_sum(reg_psum_17_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_29( .activation_in(reg_activation_17_28), .weight_in(reg_weight_16_29), .partial_sum_in(reg_psum_16_29), .reg_activation(reg_activation_17_29), .reg_weight(reg_weight_17_29), .reg_partial_sum(reg_psum_17_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_30( .activation_in(reg_activation_17_29), .weight_in(reg_weight_16_30), .partial_sum_in(reg_psum_16_30), .reg_activation(reg_activation_17_30), .reg_weight(reg_weight_17_30), .reg_partial_sum(reg_psum_17_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U17_31( .activation_in(reg_activation_17_30), .weight_in(reg_weight_16_31), .partial_sum_in(reg_psum_16_31), .reg_weight(reg_weight_17_31), .reg_partial_sum(reg_psum_17_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_0( .activation_in(in_activation_18), .weight_in(reg_weight_17_0), .partial_sum_in(reg_psum_17_0), .reg_activation(reg_activation_18_0), .reg_weight(reg_weight_18_0), .reg_partial_sum(reg_psum_18_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_1( .activation_in(reg_activation_18_0), .weight_in(reg_weight_17_1), .partial_sum_in(reg_psum_17_1), .reg_activation(reg_activation_18_1), .reg_weight(reg_weight_18_1), .reg_partial_sum(reg_psum_18_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_2( .activation_in(reg_activation_18_1), .weight_in(reg_weight_17_2), .partial_sum_in(reg_psum_17_2), .reg_activation(reg_activation_18_2), .reg_weight(reg_weight_18_2), .reg_partial_sum(reg_psum_18_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_3( .activation_in(reg_activation_18_2), .weight_in(reg_weight_17_3), .partial_sum_in(reg_psum_17_3), .reg_activation(reg_activation_18_3), .reg_weight(reg_weight_18_3), .reg_partial_sum(reg_psum_18_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_4( .activation_in(reg_activation_18_3), .weight_in(reg_weight_17_4), .partial_sum_in(reg_psum_17_4), .reg_activation(reg_activation_18_4), .reg_weight(reg_weight_18_4), .reg_partial_sum(reg_psum_18_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_5( .activation_in(reg_activation_18_4), .weight_in(reg_weight_17_5), .partial_sum_in(reg_psum_17_5), .reg_activation(reg_activation_18_5), .reg_weight(reg_weight_18_5), .reg_partial_sum(reg_psum_18_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_6( .activation_in(reg_activation_18_5), .weight_in(reg_weight_17_6), .partial_sum_in(reg_psum_17_6), .reg_activation(reg_activation_18_6), .reg_weight(reg_weight_18_6), .reg_partial_sum(reg_psum_18_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_7( .activation_in(reg_activation_18_6), .weight_in(reg_weight_17_7), .partial_sum_in(reg_psum_17_7), .reg_activation(reg_activation_18_7), .reg_weight(reg_weight_18_7), .reg_partial_sum(reg_psum_18_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_8( .activation_in(reg_activation_18_7), .weight_in(reg_weight_17_8), .partial_sum_in(reg_psum_17_8), .reg_activation(reg_activation_18_8), .reg_weight(reg_weight_18_8), .reg_partial_sum(reg_psum_18_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_9( .activation_in(reg_activation_18_8), .weight_in(reg_weight_17_9), .partial_sum_in(reg_psum_17_9), .reg_activation(reg_activation_18_9), .reg_weight(reg_weight_18_9), .reg_partial_sum(reg_psum_18_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_10( .activation_in(reg_activation_18_9), .weight_in(reg_weight_17_10), .partial_sum_in(reg_psum_17_10), .reg_activation(reg_activation_18_10), .reg_weight(reg_weight_18_10), .reg_partial_sum(reg_psum_18_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_11( .activation_in(reg_activation_18_10), .weight_in(reg_weight_17_11), .partial_sum_in(reg_psum_17_11), .reg_activation(reg_activation_18_11), .reg_weight(reg_weight_18_11), .reg_partial_sum(reg_psum_18_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_12( .activation_in(reg_activation_18_11), .weight_in(reg_weight_17_12), .partial_sum_in(reg_psum_17_12), .reg_activation(reg_activation_18_12), .reg_weight(reg_weight_18_12), .reg_partial_sum(reg_psum_18_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_13( .activation_in(reg_activation_18_12), .weight_in(reg_weight_17_13), .partial_sum_in(reg_psum_17_13), .reg_activation(reg_activation_18_13), .reg_weight(reg_weight_18_13), .reg_partial_sum(reg_psum_18_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_14( .activation_in(reg_activation_18_13), .weight_in(reg_weight_17_14), .partial_sum_in(reg_psum_17_14), .reg_activation(reg_activation_18_14), .reg_weight(reg_weight_18_14), .reg_partial_sum(reg_psum_18_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_15( .activation_in(reg_activation_18_14), .weight_in(reg_weight_17_15), .partial_sum_in(reg_psum_17_15), .reg_activation(reg_activation_18_15), .reg_weight(reg_weight_18_15), .reg_partial_sum(reg_psum_18_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_16( .activation_in(reg_activation_18_15), .weight_in(reg_weight_17_16), .partial_sum_in(reg_psum_17_16), .reg_activation(reg_activation_18_16), .reg_weight(reg_weight_18_16), .reg_partial_sum(reg_psum_18_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_17( .activation_in(reg_activation_18_16), .weight_in(reg_weight_17_17), .partial_sum_in(reg_psum_17_17), .reg_activation(reg_activation_18_17), .reg_weight(reg_weight_18_17), .reg_partial_sum(reg_psum_18_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_18( .activation_in(reg_activation_18_17), .weight_in(reg_weight_17_18), .partial_sum_in(reg_psum_17_18), .reg_activation(reg_activation_18_18), .reg_weight(reg_weight_18_18), .reg_partial_sum(reg_psum_18_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_19( .activation_in(reg_activation_18_18), .weight_in(reg_weight_17_19), .partial_sum_in(reg_psum_17_19), .reg_activation(reg_activation_18_19), .reg_weight(reg_weight_18_19), .reg_partial_sum(reg_psum_18_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_20( .activation_in(reg_activation_18_19), .weight_in(reg_weight_17_20), .partial_sum_in(reg_psum_17_20), .reg_activation(reg_activation_18_20), .reg_weight(reg_weight_18_20), .reg_partial_sum(reg_psum_18_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_21( .activation_in(reg_activation_18_20), .weight_in(reg_weight_17_21), .partial_sum_in(reg_psum_17_21), .reg_activation(reg_activation_18_21), .reg_weight(reg_weight_18_21), .reg_partial_sum(reg_psum_18_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_22( .activation_in(reg_activation_18_21), .weight_in(reg_weight_17_22), .partial_sum_in(reg_psum_17_22), .reg_activation(reg_activation_18_22), .reg_weight(reg_weight_18_22), .reg_partial_sum(reg_psum_18_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_23( .activation_in(reg_activation_18_22), .weight_in(reg_weight_17_23), .partial_sum_in(reg_psum_17_23), .reg_activation(reg_activation_18_23), .reg_weight(reg_weight_18_23), .reg_partial_sum(reg_psum_18_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_24( .activation_in(reg_activation_18_23), .weight_in(reg_weight_17_24), .partial_sum_in(reg_psum_17_24), .reg_activation(reg_activation_18_24), .reg_weight(reg_weight_18_24), .reg_partial_sum(reg_psum_18_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_25( .activation_in(reg_activation_18_24), .weight_in(reg_weight_17_25), .partial_sum_in(reg_psum_17_25), .reg_activation(reg_activation_18_25), .reg_weight(reg_weight_18_25), .reg_partial_sum(reg_psum_18_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_26( .activation_in(reg_activation_18_25), .weight_in(reg_weight_17_26), .partial_sum_in(reg_psum_17_26), .reg_activation(reg_activation_18_26), .reg_weight(reg_weight_18_26), .reg_partial_sum(reg_psum_18_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_27( .activation_in(reg_activation_18_26), .weight_in(reg_weight_17_27), .partial_sum_in(reg_psum_17_27), .reg_activation(reg_activation_18_27), .reg_weight(reg_weight_18_27), .reg_partial_sum(reg_psum_18_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_28( .activation_in(reg_activation_18_27), .weight_in(reg_weight_17_28), .partial_sum_in(reg_psum_17_28), .reg_activation(reg_activation_18_28), .reg_weight(reg_weight_18_28), .reg_partial_sum(reg_psum_18_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_29( .activation_in(reg_activation_18_28), .weight_in(reg_weight_17_29), .partial_sum_in(reg_psum_17_29), .reg_activation(reg_activation_18_29), .reg_weight(reg_weight_18_29), .reg_partial_sum(reg_psum_18_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_30( .activation_in(reg_activation_18_29), .weight_in(reg_weight_17_30), .partial_sum_in(reg_psum_17_30), .reg_activation(reg_activation_18_30), .reg_weight(reg_weight_18_30), .reg_partial_sum(reg_psum_18_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U18_31( .activation_in(reg_activation_18_30), .weight_in(reg_weight_17_31), .partial_sum_in(reg_psum_17_31), .reg_weight(reg_weight_18_31), .reg_partial_sum(reg_psum_18_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_0( .activation_in(in_activation_19), .weight_in(reg_weight_18_0), .partial_sum_in(reg_psum_18_0), .reg_activation(reg_activation_19_0), .reg_weight(reg_weight_19_0), .reg_partial_sum(reg_psum_19_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_1( .activation_in(reg_activation_19_0), .weight_in(reg_weight_18_1), .partial_sum_in(reg_psum_18_1), .reg_activation(reg_activation_19_1), .reg_weight(reg_weight_19_1), .reg_partial_sum(reg_psum_19_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_2( .activation_in(reg_activation_19_1), .weight_in(reg_weight_18_2), .partial_sum_in(reg_psum_18_2), .reg_activation(reg_activation_19_2), .reg_weight(reg_weight_19_2), .reg_partial_sum(reg_psum_19_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_3( .activation_in(reg_activation_19_2), .weight_in(reg_weight_18_3), .partial_sum_in(reg_psum_18_3), .reg_activation(reg_activation_19_3), .reg_weight(reg_weight_19_3), .reg_partial_sum(reg_psum_19_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_4( .activation_in(reg_activation_19_3), .weight_in(reg_weight_18_4), .partial_sum_in(reg_psum_18_4), .reg_activation(reg_activation_19_4), .reg_weight(reg_weight_19_4), .reg_partial_sum(reg_psum_19_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_5( .activation_in(reg_activation_19_4), .weight_in(reg_weight_18_5), .partial_sum_in(reg_psum_18_5), .reg_activation(reg_activation_19_5), .reg_weight(reg_weight_19_5), .reg_partial_sum(reg_psum_19_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_6( .activation_in(reg_activation_19_5), .weight_in(reg_weight_18_6), .partial_sum_in(reg_psum_18_6), .reg_activation(reg_activation_19_6), .reg_weight(reg_weight_19_6), .reg_partial_sum(reg_psum_19_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_7( .activation_in(reg_activation_19_6), .weight_in(reg_weight_18_7), .partial_sum_in(reg_psum_18_7), .reg_activation(reg_activation_19_7), .reg_weight(reg_weight_19_7), .reg_partial_sum(reg_psum_19_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_8( .activation_in(reg_activation_19_7), .weight_in(reg_weight_18_8), .partial_sum_in(reg_psum_18_8), .reg_activation(reg_activation_19_8), .reg_weight(reg_weight_19_8), .reg_partial_sum(reg_psum_19_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_9( .activation_in(reg_activation_19_8), .weight_in(reg_weight_18_9), .partial_sum_in(reg_psum_18_9), .reg_activation(reg_activation_19_9), .reg_weight(reg_weight_19_9), .reg_partial_sum(reg_psum_19_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_10( .activation_in(reg_activation_19_9), .weight_in(reg_weight_18_10), .partial_sum_in(reg_psum_18_10), .reg_activation(reg_activation_19_10), .reg_weight(reg_weight_19_10), .reg_partial_sum(reg_psum_19_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_11( .activation_in(reg_activation_19_10), .weight_in(reg_weight_18_11), .partial_sum_in(reg_psum_18_11), .reg_activation(reg_activation_19_11), .reg_weight(reg_weight_19_11), .reg_partial_sum(reg_psum_19_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_12( .activation_in(reg_activation_19_11), .weight_in(reg_weight_18_12), .partial_sum_in(reg_psum_18_12), .reg_activation(reg_activation_19_12), .reg_weight(reg_weight_19_12), .reg_partial_sum(reg_psum_19_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_13( .activation_in(reg_activation_19_12), .weight_in(reg_weight_18_13), .partial_sum_in(reg_psum_18_13), .reg_activation(reg_activation_19_13), .reg_weight(reg_weight_19_13), .reg_partial_sum(reg_psum_19_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_14( .activation_in(reg_activation_19_13), .weight_in(reg_weight_18_14), .partial_sum_in(reg_psum_18_14), .reg_activation(reg_activation_19_14), .reg_weight(reg_weight_19_14), .reg_partial_sum(reg_psum_19_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_15( .activation_in(reg_activation_19_14), .weight_in(reg_weight_18_15), .partial_sum_in(reg_psum_18_15), .reg_activation(reg_activation_19_15), .reg_weight(reg_weight_19_15), .reg_partial_sum(reg_psum_19_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_16( .activation_in(reg_activation_19_15), .weight_in(reg_weight_18_16), .partial_sum_in(reg_psum_18_16), .reg_activation(reg_activation_19_16), .reg_weight(reg_weight_19_16), .reg_partial_sum(reg_psum_19_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_17( .activation_in(reg_activation_19_16), .weight_in(reg_weight_18_17), .partial_sum_in(reg_psum_18_17), .reg_activation(reg_activation_19_17), .reg_weight(reg_weight_19_17), .reg_partial_sum(reg_psum_19_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_18( .activation_in(reg_activation_19_17), .weight_in(reg_weight_18_18), .partial_sum_in(reg_psum_18_18), .reg_activation(reg_activation_19_18), .reg_weight(reg_weight_19_18), .reg_partial_sum(reg_psum_19_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_19( .activation_in(reg_activation_19_18), .weight_in(reg_weight_18_19), .partial_sum_in(reg_psum_18_19), .reg_activation(reg_activation_19_19), .reg_weight(reg_weight_19_19), .reg_partial_sum(reg_psum_19_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_20( .activation_in(reg_activation_19_19), .weight_in(reg_weight_18_20), .partial_sum_in(reg_psum_18_20), .reg_activation(reg_activation_19_20), .reg_weight(reg_weight_19_20), .reg_partial_sum(reg_psum_19_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_21( .activation_in(reg_activation_19_20), .weight_in(reg_weight_18_21), .partial_sum_in(reg_psum_18_21), .reg_activation(reg_activation_19_21), .reg_weight(reg_weight_19_21), .reg_partial_sum(reg_psum_19_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_22( .activation_in(reg_activation_19_21), .weight_in(reg_weight_18_22), .partial_sum_in(reg_psum_18_22), .reg_activation(reg_activation_19_22), .reg_weight(reg_weight_19_22), .reg_partial_sum(reg_psum_19_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_23( .activation_in(reg_activation_19_22), .weight_in(reg_weight_18_23), .partial_sum_in(reg_psum_18_23), .reg_activation(reg_activation_19_23), .reg_weight(reg_weight_19_23), .reg_partial_sum(reg_psum_19_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_24( .activation_in(reg_activation_19_23), .weight_in(reg_weight_18_24), .partial_sum_in(reg_psum_18_24), .reg_activation(reg_activation_19_24), .reg_weight(reg_weight_19_24), .reg_partial_sum(reg_psum_19_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_25( .activation_in(reg_activation_19_24), .weight_in(reg_weight_18_25), .partial_sum_in(reg_psum_18_25), .reg_activation(reg_activation_19_25), .reg_weight(reg_weight_19_25), .reg_partial_sum(reg_psum_19_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_26( .activation_in(reg_activation_19_25), .weight_in(reg_weight_18_26), .partial_sum_in(reg_psum_18_26), .reg_activation(reg_activation_19_26), .reg_weight(reg_weight_19_26), .reg_partial_sum(reg_psum_19_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_27( .activation_in(reg_activation_19_26), .weight_in(reg_weight_18_27), .partial_sum_in(reg_psum_18_27), .reg_activation(reg_activation_19_27), .reg_weight(reg_weight_19_27), .reg_partial_sum(reg_psum_19_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_28( .activation_in(reg_activation_19_27), .weight_in(reg_weight_18_28), .partial_sum_in(reg_psum_18_28), .reg_activation(reg_activation_19_28), .reg_weight(reg_weight_19_28), .reg_partial_sum(reg_psum_19_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_29( .activation_in(reg_activation_19_28), .weight_in(reg_weight_18_29), .partial_sum_in(reg_psum_18_29), .reg_activation(reg_activation_19_29), .reg_weight(reg_weight_19_29), .reg_partial_sum(reg_psum_19_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_30( .activation_in(reg_activation_19_29), .weight_in(reg_weight_18_30), .partial_sum_in(reg_psum_18_30), .reg_activation(reg_activation_19_30), .reg_weight(reg_weight_19_30), .reg_partial_sum(reg_psum_19_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U19_31( .activation_in(reg_activation_19_30), .weight_in(reg_weight_18_31), .partial_sum_in(reg_psum_18_31), .reg_weight(reg_weight_19_31), .reg_partial_sum(reg_psum_19_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_0( .activation_in(in_activation_20), .weight_in(reg_weight_19_0), .partial_sum_in(fault_reg_psum_19_0), .reg_activation(reg_activation_20_0), .reg_weight(reg_weight_20_0), .reg_partial_sum(reg_psum_20_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_1( .activation_in(reg_activation_20_0), .weight_in(reg_weight_19_1), .partial_sum_in(reg_psum_19_1), .reg_activation(reg_activation_20_1), .reg_weight(reg_weight_20_1), .reg_partial_sum(reg_psum_20_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_2( .activation_in(reg_activation_20_1), .weight_in(reg_weight_19_2), .partial_sum_in(reg_psum_19_2), .reg_activation(reg_activation_20_2), .reg_weight(reg_weight_20_2), .reg_partial_sum(reg_psum_20_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_3( .activation_in(reg_activation_20_2), .weight_in(reg_weight_19_3), .partial_sum_in(reg_psum_19_3), .reg_activation(reg_activation_20_3), .reg_weight(reg_weight_20_3), .reg_partial_sum(reg_psum_20_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_4( .activation_in(reg_activation_20_3), .weight_in(reg_weight_19_4), .partial_sum_in(reg_psum_19_4), .reg_activation(reg_activation_20_4), .reg_weight(reg_weight_20_4), .reg_partial_sum(reg_psum_20_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_5( .activation_in(reg_activation_20_4), .weight_in(reg_weight_19_5), .partial_sum_in(reg_psum_19_5), .reg_activation(reg_activation_20_5), .reg_weight(reg_weight_20_5), .reg_partial_sum(reg_psum_20_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_6( .activation_in(reg_activation_20_5), .weight_in(reg_weight_19_6), .partial_sum_in(reg_psum_19_6), .reg_activation(reg_activation_20_6), .reg_weight(reg_weight_20_6), .reg_partial_sum(reg_psum_20_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_7( .activation_in(reg_activation_20_6), .weight_in(reg_weight_19_7), .partial_sum_in(reg_psum_19_7), .reg_activation(reg_activation_20_7), .reg_weight(reg_weight_20_7), .reg_partial_sum(reg_psum_20_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_8( .activation_in(reg_activation_20_7), .weight_in(reg_weight_19_8), .partial_sum_in(reg_psum_19_8), .reg_activation(reg_activation_20_8), .reg_weight(reg_weight_20_8), .reg_partial_sum(reg_psum_20_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_9( .activation_in(reg_activation_20_8), .weight_in(reg_weight_19_9), .partial_sum_in(reg_psum_19_9), .reg_activation(reg_activation_20_9), .reg_weight(reg_weight_20_9), .reg_partial_sum(reg_psum_20_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_10( .activation_in(reg_activation_20_9), .weight_in(reg_weight_19_10), .partial_sum_in(reg_psum_19_10), .reg_activation(reg_activation_20_10), .reg_weight(reg_weight_20_10), .reg_partial_sum(reg_psum_20_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_11( .activation_in(reg_activation_20_10), .weight_in(reg_weight_19_11), .partial_sum_in(reg_psum_19_11), .reg_activation(reg_activation_20_11), .reg_weight(reg_weight_20_11), .reg_partial_sum(reg_psum_20_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_12( .activation_in(reg_activation_20_11), .weight_in(reg_weight_19_12), .partial_sum_in(reg_psum_19_12), .reg_activation(reg_activation_20_12), .reg_weight(reg_weight_20_12), .reg_partial_sum(reg_psum_20_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_13( .activation_in(reg_activation_20_12), .weight_in(reg_weight_19_13), .partial_sum_in(reg_psum_19_13), .reg_activation(reg_activation_20_13), .reg_weight(reg_weight_20_13), .reg_partial_sum(reg_psum_20_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_14( .activation_in(reg_activation_20_13), .weight_in(reg_weight_19_14), .partial_sum_in(reg_psum_19_14), .reg_activation(reg_activation_20_14), .reg_weight(reg_weight_20_14), .reg_partial_sum(reg_psum_20_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_15( .activation_in(reg_activation_20_14), .weight_in(reg_weight_19_15), .partial_sum_in(reg_psum_19_15), .reg_activation(reg_activation_20_15), .reg_weight(reg_weight_20_15), .reg_partial_sum(reg_psum_20_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_16( .activation_in(reg_activation_20_15), .weight_in(reg_weight_19_16), .partial_sum_in(reg_psum_19_16), .reg_activation(reg_activation_20_16), .reg_weight(reg_weight_20_16), .reg_partial_sum(reg_psum_20_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_17( .activation_in(reg_activation_20_16), .weight_in(reg_weight_19_17), .partial_sum_in(reg_psum_19_17), .reg_activation(reg_activation_20_17), .reg_weight(reg_weight_20_17), .reg_partial_sum(reg_psum_20_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_18( .activation_in(reg_activation_20_17), .weight_in(reg_weight_19_18), .partial_sum_in(reg_psum_19_18), .reg_activation(reg_activation_20_18), .reg_weight(reg_weight_20_18), .reg_partial_sum(reg_psum_20_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_19( .activation_in(reg_activation_20_18), .weight_in(reg_weight_19_19), .partial_sum_in(reg_psum_19_19), .reg_activation(reg_activation_20_19), .reg_weight(reg_weight_20_19), .reg_partial_sum(reg_psum_20_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_20( .activation_in(reg_activation_20_19), .weight_in(reg_weight_19_20), .partial_sum_in(reg_psum_19_20), .reg_activation(reg_activation_20_20), .reg_weight(reg_weight_20_20), .reg_partial_sum(reg_psum_20_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_21( .activation_in(reg_activation_20_20), .weight_in(reg_weight_19_21), .partial_sum_in(reg_psum_19_21), .reg_activation(reg_activation_20_21), .reg_weight(reg_weight_20_21), .reg_partial_sum(reg_psum_20_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_22( .activation_in(reg_activation_20_21), .weight_in(reg_weight_19_22), .partial_sum_in(reg_psum_19_22), .reg_activation(reg_activation_20_22), .reg_weight(reg_weight_20_22), .reg_partial_sum(reg_psum_20_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_23( .activation_in(reg_activation_20_22), .weight_in(reg_weight_19_23), .partial_sum_in(reg_psum_19_23), .reg_activation(reg_activation_20_23), .reg_weight(reg_weight_20_23), .reg_partial_sum(reg_psum_20_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_24( .activation_in(reg_activation_20_23), .weight_in(reg_weight_19_24), .partial_sum_in(reg_psum_19_24), .reg_activation(reg_activation_20_24), .reg_weight(reg_weight_20_24), .reg_partial_sum(reg_psum_20_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_25( .activation_in(reg_activation_20_24), .weight_in(reg_weight_19_25), .partial_sum_in(reg_psum_19_25), .reg_activation(reg_activation_20_25), .reg_weight(reg_weight_20_25), .reg_partial_sum(reg_psum_20_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_26( .activation_in(reg_activation_20_25), .weight_in(reg_weight_19_26), .partial_sum_in(reg_psum_19_26), .reg_activation(reg_activation_20_26), .reg_weight(reg_weight_20_26), .reg_partial_sum(reg_psum_20_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_27( .activation_in(reg_activation_20_26), .weight_in(reg_weight_19_27), .partial_sum_in(reg_psum_19_27), .reg_activation(reg_activation_20_27), .reg_weight(reg_weight_20_27), .reg_partial_sum(reg_psum_20_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_28( .activation_in(reg_activation_20_27), .weight_in(reg_weight_19_28), .partial_sum_in(reg_psum_19_28), .reg_activation(reg_activation_20_28), .reg_weight(reg_weight_20_28), .reg_partial_sum(reg_psum_20_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_29( .activation_in(reg_activation_20_28), .weight_in(reg_weight_19_29), .partial_sum_in(reg_psum_19_29), .reg_activation(reg_activation_20_29), .reg_weight(reg_weight_20_29), .reg_partial_sum(reg_psum_20_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_30( .activation_in(reg_activation_20_29), .weight_in(reg_weight_19_30), .partial_sum_in(reg_psum_19_30), .reg_activation(reg_activation_20_30), .reg_weight(reg_weight_20_30), .reg_partial_sum(reg_psum_20_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U20_31( .activation_in(reg_activation_20_30), .weight_in(reg_weight_19_31), .partial_sum_in(reg_psum_19_31), .reg_weight(reg_weight_20_31), .reg_partial_sum(reg_psum_20_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_0( .activation_in(in_activation_21), .weight_in(reg_weight_20_0), .partial_sum_in(reg_psum_20_0), .reg_activation(reg_activation_21_0), .reg_weight(reg_weight_21_0), .reg_partial_sum(reg_psum_21_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_1( .activation_in(reg_activation_21_0), .weight_in(reg_weight_20_1), .partial_sum_in(reg_psum_20_1), .reg_activation(reg_activation_21_1), .reg_weight(reg_weight_21_1), .reg_partial_sum(reg_psum_21_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_2( .activation_in(reg_activation_21_1), .weight_in(reg_weight_20_2), .partial_sum_in(reg_psum_20_2), .reg_activation(reg_activation_21_2), .reg_weight(reg_weight_21_2), .reg_partial_sum(reg_psum_21_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_3( .activation_in(reg_activation_21_2), .weight_in(reg_weight_20_3), .partial_sum_in(reg_psum_20_3), .reg_activation(reg_activation_21_3), .reg_weight(reg_weight_21_3), .reg_partial_sum(reg_psum_21_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_4( .activation_in(reg_activation_21_3), .weight_in(reg_weight_20_4), .partial_sum_in(reg_psum_20_4), .reg_activation(reg_activation_21_4), .reg_weight(reg_weight_21_4), .reg_partial_sum(reg_psum_21_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_5( .activation_in(reg_activation_21_4), .weight_in(reg_weight_20_5), .partial_sum_in(reg_psum_20_5), .reg_activation(reg_activation_21_5), .reg_weight(reg_weight_21_5), .reg_partial_sum(reg_psum_21_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_6( .activation_in(reg_activation_21_5), .weight_in(reg_weight_20_6), .partial_sum_in(reg_psum_20_6), .reg_activation(reg_activation_21_6), .reg_weight(reg_weight_21_6), .reg_partial_sum(reg_psum_21_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_7( .activation_in(reg_activation_21_6), .weight_in(reg_weight_20_7), .partial_sum_in(reg_psum_20_7), .reg_activation(reg_activation_21_7), .reg_weight(reg_weight_21_7), .reg_partial_sum(reg_psum_21_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_8( .activation_in(reg_activation_21_7), .weight_in(reg_weight_20_8), .partial_sum_in(reg_psum_20_8), .reg_activation(reg_activation_21_8), .reg_weight(reg_weight_21_8), .reg_partial_sum(reg_psum_21_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_9( .activation_in(reg_activation_21_8), .weight_in(reg_weight_20_9), .partial_sum_in(reg_psum_20_9), .reg_activation(reg_activation_21_9), .reg_weight(reg_weight_21_9), .reg_partial_sum(reg_psum_21_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_10( .activation_in(reg_activation_21_9), .weight_in(reg_weight_20_10), .partial_sum_in(reg_psum_20_10), .reg_activation(reg_activation_21_10), .reg_weight(reg_weight_21_10), .reg_partial_sum(reg_psum_21_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_11( .activation_in(reg_activation_21_10), .weight_in(reg_weight_20_11), .partial_sum_in(fault_reg_psum_20_11), .reg_activation(reg_activation_21_11), .reg_weight(reg_weight_21_11), .reg_partial_sum(reg_psum_21_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_12( .activation_in(reg_activation_21_11), .weight_in(reg_weight_20_12), .partial_sum_in(reg_psum_20_12), .reg_activation(reg_activation_21_12), .reg_weight(reg_weight_21_12), .reg_partial_sum(reg_psum_21_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_13( .activation_in(reg_activation_21_12), .weight_in(reg_weight_20_13), .partial_sum_in(reg_psum_20_13), .reg_activation(reg_activation_21_13), .reg_weight(reg_weight_21_13), .reg_partial_sum(reg_psum_21_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_14( .activation_in(reg_activation_21_13), .weight_in(reg_weight_20_14), .partial_sum_in(reg_psum_20_14), .reg_activation(reg_activation_21_14), .reg_weight(reg_weight_21_14), .reg_partial_sum(reg_psum_21_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_15( .activation_in(reg_activation_21_14), .weight_in(reg_weight_20_15), .partial_sum_in(reg_psum_20_15), .reg_activation(reg_activation_21_15), .reg_weight(reg_weight_21_15), .reg_partial_sum(reg_psum_21_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_16( .activation_in(reg_activation_21_15), .weight_in(reg_weight_20_16), .partial_sum_in(reg_psum_20_16), .reg_activation(reg_activation_21_16), .reg_weight(reg_weight_21_16), .reg_partial_sum(reg_psum_21_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_17( .activation_in(reg_activation_21_16), .weight_in(reg_weight_20_17), .partial_sum_in(reg_psum_20_17), .reg_activation(reg_activation_21_17), .reg_weight(reg_weight_21_17), .reg_partial_sum(reg_psum_21_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_18( .activation_in(reg_activation_21_17), .weight_in(reg_weight_20_18), .partial_sum_in(reg_psum_20_18), .reg_activation(reg_activation_21_18), .reg_weight(reg_weight_21_18), .reg_partial_sum(reg_psum_21_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_19( .activation_in(reg_activation_21_18), .weight_in(reg_weight_20_19), .partial_sum_in(reg_psum_20_19), .reg_activation(reg_activation_21_19), .reg_weight(reg_weight_21_19), .reg_partial_sum(reg_psum_21_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_20( .activation_in(reg_activation_21_19), .weight_in(reg_weight_20_20), .partial_sum_in(reg_psum_20_20), .reg_activation(reg_activation_21_20), .reg_weight(reg_weight_21_20), .reg_partial_sum(reg_psum_21_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_21( .activation_in(reg_activation_21_20), .weight_in(reg_weight_20_21), .partial_sum_in(reg_psum_20_21), .reg_activation(reg_activation_21_21), .reg_weight(reg_weight_21_21), .reg_partial_sum(reg_psum_21_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_22( .activation_in(reg_activation_21_21), .weight_in(reg_weight_20_22), .partial_sum_in(reg_psum_20_22), .reg_activation(reg_activation_21_22), .reg_weight(reg_weight_21_22), .reg_partial_sum(reg_psum_21_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_23( .activation_in(reg_activation_21_22), .weight_in(reg_weight_20_23), .partial_sum_in(reg_psum_20_23), .reg_activation(reg_activation_21_23), .reg_weight(reg_weight_21_23), .reg_partial_sum(reg_psum_21_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_24( .activation_in(reg_activation_21_23), .weight_in(reg_weight_20_24), .partial_sum_in(reg_psum_20_24), .reg_activation(reg_activation_21_24), .reg_weight(reg_weight_21_24), .reg_partial_sum(reg_psum_21_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_25( .activation_in(reg_activation_21_24), .weight_in(reg_weight_20_25), .partial_sum_in(reg_psum_20_25), .reg_activation(reg_activation_21_25), .reg_weight(reg_weight_21_25), .reg_partial_sum(reg_psum_21_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_26( .activation_in(reg_activation_21_25), .weight_in(reg_weight_20_26), .partial_sum_in(reg_psum_20_26), .reg_activation(reg_activation_21_26), .reg_weight(reg_weight_21_26), .reg_partial_sum(reg_psum_21_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_27( .activation_in(reg_activation_21_26), .weight_in(reg_weight_20_27), .partial_sum_in(reg_psum_20_27), .reg_activation(reg_activation_21_27), .reg_weight(reg_weight_21_27), .reg_partial_sum(reg_psum_21_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_28( .activation_in(reg_activation_21_27), .weight_in(reg_weight_20_28), .partial_sum_in(reg_psum_20_28), .reg_activation(reg_activation_21_28), .reg_weight(reg_weight_21_28), .reg_partial_sum(reg_psum_21_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_29( .activation_in(reg_activation_21_28), .weight_in(reg_weight_20_29), .partial_sum_in(reg_psum_20_29), .reg_activation(reg_activation_21_29), .reg_weight(reg_weight_21_29), .reg_partial_sum(reg_psum_21_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_30( .activation_in(reg_activation_21_29), .weight_in(reg_weight_20_30), .partial_sum_in(reg_psum_20_30), .reg_activation(reg_activation_21_30), .reg_weight(reg_weight_21_30), .reg_partial_sum(reg_psum_21_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U21_31( .activation_in(reg_activation_21_30), .weight_in(reg_weight_20_31), .partial_sum_in(reg_psum_20_31), .reg_weight(reg_weight_21_31), .reg_partial_sum(reg_psum_21_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_0( .activation_in(in_activation_22), .weight_in(reg_weight_21_0), .partial_sum_in(reg_psum_21_0), .reg_activation(reg_activation_22_0), .reg_weight(reg_weight_22_0), .reg_partial_sum(reg_psum_22_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_1( .activation_in(reg_activation_22_0), .weight_in(reg_weight_21_1), .partial_sum_in(reg_psum_21_1), .reg_activation(reg_activation_22_1), .reg_weight(reg_weight_22_1), .reg_partial_sum(reg_psum_22_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_2( .activation_in(reg_activation_22_1), .weight_in(reg_weight_21_2), .partial_sum_in(reg_psum_21_2), .reg_activation(reg_activation_22_2), .reg_weight(reg_weight_22_2), .reg_partial_sum(reg_psum_22_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_3( .activation_in(reg_activation_22_2), .weight_in(reg_weight_21_3), .partial_sum_in(reg_psum_21_3), .reg_activation(reg_activation_22_3), .reg_weight(reg_weight_22_3), .reg_partial_sum(reg_psum_22_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_4( .activation_in(reg_activation_22_3), .weight_in(reg_weight_21_4), .partial_sum_in(reg_psum_21_4), .reg_activation(reg_activation_22_4), .reg_weight(reg_weight_22_4), .reg_partial_sum(reg_psum_22_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_5( .activation_in(reg_activation_22_4), .weight_in(reg_weight_21_5), .partial_sum_in(reg_psum_21_5), .reg_activation(reg_activation_22_5), .reg_weight(reg_weight_22_5), .reg_partial_sum(reg_psum_22_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_6( .activation_in(reg_activation_22_5), .weight_in(reg_weight_21_6), .partial_sum_in(reg_psum_21_6), .reg_activation(reg_activation_22_6), .reg_weight(reg_weight_22_6), .reg_partial_sum(reg_psum_22_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_7( .activation_in(reg_activation_22_6), .weight_in(reg_weight_21_7), .partial_sum_in(reg_psum_21_7), .reg_activation(reg_activation_22_7), .reg_weight(reg_weight_22_7), .reg_partial_sum(reg_psum_22_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_8( .activation_in(reg_activation_22_7), .weight_in(reg_weight_21_8), .partial_sum_in(reg_psum_21_8), .reg_activation(reg_activation_22_8), .reg_weight(reg_weight_22_8), .reg_partial_sum(reg_psum_22_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_9( .activation_in(reg_activation_22_8), .weight_in(reg_weight_21_9), .partial_sum_in(reg_psum_21_9), .reg_activation(reg_activation_22_9), .reg_weight(reg_weight_22_9), .reg_partial_sum(reg_psum_22_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_10( .activation_in(reg_activation_22_9), .weight_in(reg_weight_21_10), .partial_sum_in(reg_psum_21_10), .reg_activation(reg_activation_22_10), .reg_weight(reg_weight_22_10), .reg_partial_sum(reg_psum_22_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_11( .activation_in(reg_activation_22_10), .weight_in(reg_weight_21_11), .partial_sum_in(reg_psum_21_11), .reg_activation(reg_activation_22_11), .reg_weight(reg_weight_22_11), .reg_partial_sum(reg_psum_22_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_12( .activation_in(reg_activation_22_11), .weight_in(reg_weight_21_12), .partial_sum_in(reg_psum_21_12), .reg_activation(reg_activation_22_12), .reg_weight(reg_weight_22_12), .reg_partial_sum(reg_psum_22_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_13( .activation_in(reg_activation_22_12), .weight_in(reg_weight_21_13), .partial_sum_in(reg_psum_21_13), .reg_activation(reg_activation_22_13), .reg_weight(reg_weight_22_13), .reg_partial_sum(reg_psum_22_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_14( .activation_in(reg_activation_22_13), .weight_in(reg_weight_21_14), .partial_sum_in(reg_psum_21_14), .reg_activation(reg_activation_22_14), .reg_weight(reg_weight_22_14), .reg_partial_sum(reg_psum_22_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_15( .activation_in(reg_activation_22_14), .weight_in(reg_weight_21_15), .partial_sum_in(reg_psum_21_15), .reg_activation(reg_activation_22_15), .reg_weight(reg_weight_22_15), .reg_partial_sum(reg_psum_22_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_16( .activation_in(reg_activation_22_15), .weight_in(reg_weight_21_16), .partial_sum_in(reg_psum_21_16), .reg_activation(reg_activation_22_16), .reg_weight(reg_weight_22_16), .reg_partial_sum(reg_psum_22_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_17( .activation_in(reg_activation_22_16), .weight_in(reg_weight_21_17), .partial_sum_in(fault_reg_psum_21_17), .reg_activation(reg_activation_22_17), .reg_weight(reg_weight_22_17), .reg_partial_sum(reg_psum_22_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_18( .activation_in(reg_activation_22_17), .weight_in(reg_weight_21_18), .partial_sum_in(reg_psum_21_18), .reg_activation(reg_activation_22_18), .reg_weight(reg_weight_22_18), .reg_partial_sum(reg_psum_22_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_19( .activation_in(reg_activation_22_18), .weight_in(reg_weight_21_19), .partial_sum_in(reg_psum_21_19), .reg_activation(reg_activation_22_19), .reg_weight(reg_weight_22_19), .reg_partial_sum(reg_psum_22_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_20( .activation_in(reg_activation_22_19), .weight_in(reg_weight_21_20), .partial_sum_in(reg_psum_21_20), .reg_activation(reg_activation_22_20), .reg_weight(reg_weight_22_20), .reg_partial_sum(reg_psum_22_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_21( .activation_in(reg_activation_22_20), .weight_in(reg_weight_21_21), .partial_sum_in(reg_psum_21_21), .reg_activation(reg_activation_22_21), .reg_weight(reg_weight_22_21), .reg_partial_sum(reg_psum_22_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_22( .activation_in(reg_activation_22_21), .weight_in(reg_weight_21_22), .partial_sum_in(reg_psum_21_22), .reg_activation(reg_activation_22_22), .reg_weight(reg_weight_22_22), .reg_partial_sum(reg_psum_22_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_23( .activation_in(reg_activation_22_22), .weight_in(reg_weight_21_23), .partial_sum_in(reg_psum_21_23), .reg_activation(reg_activation_22_23), .reg_weight(reg_weight_22_23), .reg_partial_sum(reg_psum_22_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_24( .activation_in(reg_activation_22_23), .weight_in(reg_weight_21_24), .partial_sum_in(reg_psum_21_24), .reg_activation(reg_activation_22_24), .reg_weight(reg_weight_22_24), .reg_partial_sum(reg_psum_22_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_25( .activation_in(reg_activation_22_24), .weight_in(reg_weight_21_25), .partial_sum_in(reg_psum_21_25), .reg_activation(reg_activation_22_25), .reg_weight(reg_weight_22_25), .reg_partial_sum(reg_psum_22_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_26( .activation_in(reg_activation_22_25), .weight_in(reg_weight_21_26), .partial_sum_in(reg_psum_21_26), .reg_activation(reg_activation_22_26), .reg_weight(reg_weight_22_26), .reg_partial_sum(reg_psum_22_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_27( .activation_in(reg_activation_22_26), .weight_in(reg_weight_21_27), .partial_sum_in(reg_psum_21_27), .reg_activation(reg_activation_22_27), .reg_weight(reg_weight_22_27), .reg_partial_sum(reg_psum_22_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_28( .activation_in(reg_activation_22_27), .weight_in(reg_weight_21_28), .partial_sum_in(reg_psum_21_28), .reg_activation(reg_activation_22_28), .reg_weight(reg_weight_22_28), .reg_partial_sum(reg_psum_22_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_29( .activation_in(reg_activation_22_28), .weight_in(reg_weight_21_29), .partial_sum_in(reg_psum_21_29), .reg_activation(reg_activation_22_29), .reg_weight(reg_weight_22_29), .reg_partial_sum(reg_psum_22_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_30( .activation_in(reg_activation_22_29), .weight_in(reg_weight_21_30), .partial_sum_in(fault_reg_psum_21_30), .reg_activation(reg_activation_22_30), .reg_weight(reg_weight_22_30), .reg_partial_sum(reg_psum_22_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U22_31( .activation_in(reg_activation_22_30), .weight_in(reg_weight_21_31), .partial_sum_in(reg_psum_21_31), .reg_weight(reg_weight_22_31), .reg_partial_sum(reg_psum_22_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_0( .activation_in(in_activation_23), .weight_in(reg_weight_22_0), .partial_sum_in(reg_psum_22_0), .reg_activation(reg_activation_23_0), .reg_weight(reg_weight_23_0), .reg_partial_sum(reg_psum_23_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_1( .activation_in(reg_activation_23_0), .weight_in(reg_weight_22_1), .partial_sum_in(reg_psum_22_1), .reg_activation(reg_activation_23_1), .reg_weight(reg_weight_23_1), .reg_partial_sum(reg_psum_23_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_2( .activation_in(reg_activation_23_1), .weight_in(reg_weight_22_2), .partial_sum_in(reg_psum_22_2), .reg_activation(reg_activation_23_2), .reg_weight(reg_weight_23_2), .reg_partial_sum(reg_psum_23_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_3( .activation_in(reg_activation_23_2), .weight_in(reg_weight_22_3), .partial_sum_in(reg_psum_22_3), .reg_activation(reg_activation_23_3), .reg_weight(reg_weight_23_3), .reg_partial_sum(reg_psum_23_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_4( .activation_in(reg_activation_23_3), .weight_in(reg_weight_22_4), .partial_sum_in(reg_psum_22_4), .reg_activation(reg_activation_23_4), .reg_weight(reg_weight_23_4), .reg_partial_sum(reg_psum_23_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_5( .activation_in(reg_activation_23_4), .weight_in(reg_weight_22_5), .partial_sum_in(reg_psum_22_5), .reg_activation(reg_activation_23_5), .reg_weight(reg_weight_23_5), .reg_partial_sum(reg_psum_23_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_6( .activation_in(reg_activation_23_5), .weight_in(reg_weight_22_6), .partial_sum_in(reg_psum_22_6), .reg_activation(reg_activation_23_6), .reg_weight(reg_weight_23_6), .reg_partial_sum(reg_psum_23_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_7( .activation_in(reg_activation_23_6), .weight_in(reg_weight_22_7), .partial_sum_in(reg_psum_22_7), .reg_activation(reg_activation_23_7), .reg_weight(reg_weight_23_7), .reg_partial_sum(reg_psum_23_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_8( .activation_in(reg_activation_23_7), .weight_in(reg_weight_22_8), .partial_sum_in(reg_psum_22_8), .reg_activation(reg_activation_23_8), .reg_weight(reg_weight_23_8), .reg_partial_sum(reg_psum_23_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_9( .activation_in(reg_activation_23_8), .weight_in(reg_weight_22_9), .partial_sum_in(reg_psum_22_9), .reg_activation(reg_activation_23_9), .reg_weight(reg_weight_23_9), .reg_partial_sum(reg_psum_23_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_10( .activation_in(reg_activation_23_9), .weight_in(reg_weight_22_10), .partial_sum_in(reg_psum_22_10), .reg_activation(reg_activation_23_10), .reg_weight(reg_weight_23_10), .reg_partial_sum(reg_psum_23_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_11( .activation_in(reg_activation_23_10), .weight_in(reg_weight_22_11), .partial_sum_in(reg_psum_22_11), .reg_activation(reg_activation_23_11), .reg_weight(reg_weight_23_11), .reg_partial_sum(reg_psum_23_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_12( .activation_in(reg_activation_23_11), .weight_in(reg_weight_22_12), .partial_sum_in(reg_psum_22_12), .reg_activation(reg_activation_23_12), .reg_weight(reg_weight_23_12), .reg_partial_sum(reg_psum_23_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_13( .activation_in(reg_activation_23_12), .weight_in(reg_weight_22_13), .partial_sum_in(reg_psum_22_13), .reg_activation(reg_activation_23_13), .reg_weight(reg_weight_23_13), .reg_partial_sum(reg_psum_23_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_14( .activation_in(reg_activation_23_13), .weight_in(reg_weight_22_14), .partial_sum_in(reg_psum_22_14), .reg_activation(reg_activation_23_14), .reg_weight(reg_weight_23_14), .reg_partial_sum(reg_psum_23_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_15( .activation_in(reg_activation_23_14), .weight_in(reg_weight_22_15), .partial_sum_in(reg_psum_22_15), .reg_activation(reg_activation_23_15), .reg_weight(reg_weight_23_15), .reg_partial_sum(reg_psum_23_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_16( .activation_in(reg_activation_23_15), .weight_in(reg_weight_22_16), .partial_sum_in(reg_psum_22_16), .reg_activation(reg_activation_23_16), .reg_weight(reg_weight_23_16), .reg_partial_sum(reg_psum_23_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_17( .activation_in(reg_activation_23_16), .weight_in(reg_weight_22_17), .partial_sum_in(reg_psum_22_17), .reg_activation(reg_activation_23_17), .reg_weight(reg_weight_23_17), .reg_partial_sum(reg_psum_23_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_18( .activation_in(reg_activation_23_17), .weight_in(reg_weight_22_18), .partial_sum_in(reg_psum_22_18), .reg_activation(reg_activation_23_18), .reg_weight(reg_weight_23_18), .reg_partial_sum(reg_psum_23_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_19( .activation_in(reg_activation_23_18), .weight_in(reg_weight_22_19), .partial_sum_in(reg_psum_22_19), .reg_activation(reg_activation_23_19), .reg_weight(reg_weight_23_19), .reg_partial_sum(reg_psum_23_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_20( .activation_in(reg_activation_23_19), .weight_in(reg_weight_22_20), .partial_sum_in(reg_psum_22_20), .reg_activation(reg_activation_23_20), .reg_weight(reg_weight_23_20), .reg_partial_sum(reg_psum_23_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_21( .activation_in(reg_activation_23_20), .weight_in(reg_weight_22_21), .partial_sum_in(reg_psum_22_21), .reg_activation(reg_activation_23_21), .reg_weight(reg_weight_23_21), .reg_partial_sum(reg_psum_23_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_22( .activation_in(reg_activation_23_21), .weight_in(reg_weight_22_22), .partial_sum_in(reg_psum_22_22), .reg_activation(reg_activation_23_22), .reg_weight(reg_weight_23_22), .reg_partial_sum(reg_psum_23_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_23( .activation_in(reg_activation_23_22), .weight_in(reg_weight_22_23), .partial_sum_in(reg_psum_22_23), .reg_activation(reg_activation_23_23), .reg_weight(reg_weight_23_23), .reg_partial_sum(reg_psum_23_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_24( .activation_in(reg_activation_23_23), .weight_in(reg_weight_22_24), .partial_sum_in(reg_psum_22_24), .reg_activation(reg_activation_23_24), .reg_weight(reg_weight_23_24), .reg_partial_sum(reg_psum_23_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_25( .activation_in(reg_activation_23_24), .weight_in(reg_weight_22_25), .partial_sum_in(reg_psum_22_25), .reg_activation(reg_activation_23_25), .reg_weight(reg_weight_23_25), .reg_partial_sum(reg_psum_23_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_26( .activation_in(reg_activation_23_25), .weight_in(reg_weight_22_26), .partial_sum_in(reg_psum_22_26), .reg_activation(reg_activation_23_26), .reg_weight(reg_weight_23_26), .reg_partial_sum(reg_psum_23_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_27( .activation_in(reg_activation_23_26), .weight_in(reg_weight_22_27), .partial_sum_in(reg_psum_22_27), .reg_activation(reg_activation_23_27), .reg_weight(reg_weight_23_27), .reg_partial_sum(reg_psum_23_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_28( .activation_in(reg_activation_23_27), .weight_in(reg_weight_22_28), .partial_sum_in(reg_psum_22_28), .reg_activation(reg_activation_23_28), .reg_weight(reg_weight_23_28), .reg_partial_sum(reg_psum_23_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_29( .activation_in(reg_activation_23_28), .weight_in(reg_weight_22_29), .partial_sum_in(reg_psum_22_29), .reg_activation(reg_activation_23_29), .reg_weight(reg_weight_23_29), .reg_partial_sum(reg_psum_23_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_30( .activation_in(reg_activation_23_29), .weight_in(reg_weight_22_30), .partial_sum_in(fault_reg_psum_22_30), .reg_activation(reg_activation_23_30), .reg_weight(reg_weight_23_30), .reg_partial_sum(reg_psum_23_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U23_31( .activation_in(reg_activation_23_30), .weight_in(reg_weight_22_31), .partial_sum_in(reg_psum_22_31), .reg_weight(reg_weight_23_31), .reg_partial_sum(reg_psum_23_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_0( .activation_in(in_activation_24), .weight_in(reg_weight_23_0), .partial_sum_in(reg_psum_23_0), .reg_activation(reg_activation_24_0), .reg_weight(reg_weight_24_0), .reg_partial_sum(reg_psum_24_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_1( .activation_in(reg_activation_24_0), .weight_in(reg_weight_23_1), .partial_sum_in(reg_psum_23_1), .reg_activation(reg_activation_24_1), .reg_weight(reg_weight_24_1), .reg_partial_sum(reg_psum_24_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_2( .activation_in(reg_activation_24_1), .weight_in(reg_weight_23_2), .partial_sum_in(reg_psum_23_2), .reg_activation(reg_activation_24_2), .reg_weight(reg_weight_24_2), .reg_partial_sum(reg_psum_24_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_3( .activation_in(reg_activation_24_2), .weight_in(reg_weight_23_3), .partial_sum_in(reg_psum_23_3), .reg_activation(reg_activation_24_3), .reg_weight(reg_weight_24_3), .reg_partial_sum(reg_psum_24_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_4( .activation_in(reg_activation_24_3), .weight_in(reg_weight_23_4), .partial_sum_in(reg_psum_23_4), .reg_activation(reg_activation_24_4), .reg_weight(reg_weight_24_4), .reg_partial_sum(reg_psum_24_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_5( .activation_in(reg_activation_24_4), .weight_in(reg_weight_23_5), .partial_sum_in(reg_psum_23_5), .reg_activation(reg_activation_24_5), .reg_weight(reg_weight_24_5), .reg_partial_sum(reg_psum_24_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_6( .activation_in(reg_activation_24_5), .weight_in(reg_weight_23_6), .partial_sum_in(reg_psum_23_6), .reg_activation(reg_activation_24_6), .reg_weight(reg_weight_24_6), .reg_partial_sum(reg_psum_24_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_7( .activation_in(reg_activation_24_6), .weight_in(reg_weight_23_7), .partial_sum_in(reg_psum_23_7), .reg_activation(reg_activation_24_7), .reg_weight(reg_weight_24_7), .reg_partial_sum(reg_psum_24_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_8( .activation_in(reg_activation_24_7), .weight_in(reg_weight_23_8), .partial_sum_in(reg_psum_23_8), .reg_activation(reg_activation_24_8), .reg_weight(reg_weight_24_8), .reg_partial_sum(reg_psum_24_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_9( .activation_in(reg_activation_24_8), .weight_in(reg_weight_23_9), .partial_sum_in(reg_psum_23_9), .reg_activation(reg_activation_24_9), .reg_weight(reg_weight_24_9), .reg_partial_sum(reg_psum_24_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_10( .activation_in(reg_activation_24_9), .weight_in(reg_weight_23_10), .partial_sum_in(reg_psum_23_10), .reg_activation(reg_activation_24_10), .reg_weight(reg_weight_24_10), .reg_partial_sum(reg_psum_24_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_11( .activation_in(reg_activation_24_10), .weight_in(reg_weight_23_11), .partial_sum_in(reg_psum_23_11), .reg_activation(reg_activation_24_11), .reg_weight(reg_weight_24_11), .reg_partial_sum(reg_psum_24_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_12( .activation_in(reg_activation_24_11), .weight_in(reg_weight_23_12), .partial_sum_in(reg_psum_23_12), .reg_activation(reg_activation_24_12), .reg_weight(reg_weight_24_12), .reg_partial_sum(reg_psum_24_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_13( .activation_in(reg_activation_24_12), .weight_in(reg_weight_23_13), .partial_sum_in(reg_psum_23_13), .reg_activation(reg_activation_24_13), .reg_weight(reg_weight_24_13), .reg_partial_sum(reg_psum_24_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_14( .activation_in(reg_activation_24_13), .weight_in(reg_weight_23_14), .partial_sum_in(reg_psum_23_14), .reg_activation(reg_activation_24_14), .reg_weight(reg_weight_24_14), .reg_partial_sum(reg_psum_24_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_15( .activation_in(reg_activation_24_14), .weight_in(reg_weight_23_15), .partial_sum_in(reg_psum_23_15), .reg_activation(reg_activation_24_15), .reg_weight(reg_weight_24_15), .reg_partial_sum(reg_psum_24_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_16( .activation_in(reg_activation_24_15), .weight_in(reg_weight_23_16), .partial_sum_in(reg_psum_23_16), .reg_activation(reg_activation_24_16), .reg_weight(reg_weight_24_16), .reg_partial_sum(reg_psum_24_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_17( .activation_in(reg_activation_24_16), .weight_in(reg_weight_23_17), .partial_sum_in(reg_psum_23_17), .reg_activation(reg_activation_24_17), .reg_weight(reg_weight_24_17), .reg_partial_sum(reg_psum_24_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_18( .activation_in(reg_activation_24_17), .weight_in(reg_weight_23_18), .partial_sum_in(reg_psum_23_18), .reg_activation(reg_activation_24_18), .reg_weight(reg_weight_24_18), .reg_partial_sum(reg_psum_24_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_19( .activation_in(reg_activation_24_18), .weight_in(reg_weight_23_19), .partial_sum_in(reg_psum_23_19), .reg_activation(reg_activation_24_19), .reg_weight(reg_weight_24_19), .reg_partial_sum(reg_psum_24_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_20( .activation_in(reg_activation_24_19), .weight_in(reg_weight_23_20), .partial_sum_in(reg_psum_23_20), .reg_activation(reg_activation_24_20), .reg_weight(reg_weight_24_20), .reg_partial_sum(reg_psum_24_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_21( .activation_in(reg_activation_24_20), .weight_in(reg_weight_23_21), .partial_sum_in(reg_psum_23_21), .reg_activation(reg_activation_24_21), .reg_weight(reg_weight_24_21), .reg_partial_sum(reg_psum_24_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_22( .activation_in(reg_activation_24_21), .weight_in(reg_weight_23_22), .partial_sum_in(reg_psum_23_22), .reg_activation(reg_activation_24_22), .reg_weight(reg_weight_24_22), .reg_partial_sum(reg_psum_24_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_23( .activation_in(reg_activation_24_22), .weight_in(reg_weight_23_23), .partial_sum_in(reg_psum_23_23), .reg_activation(reg_activation_24_23), .reg_weight(reg_weight_24_23), .reg_partial_sum(reg_psum_24_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_24( .activation_in(reg_activation_24_23), .weight_in(reg_weight_23_24), .partial_sum_in(reg_psum_23_24), .reg_activation(reg_activation_24_24), .reg_weight(reg_weight_24_24), .reg_partial_sum(reg_psum_24_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_25( .activation_in(reg_activation_24_24), .weight_in(reg_weight_23_25), .partial_sum_in(reg_psum_23_25), .reg_activation(reg_activation_24_25), .reg_weight(reg_weight_24_25), .reg_partial_sum(reg_psum_24_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_26( .activation_in(reg_activation_24_25), .weight_in(reg_weight_23_26), .partial_sum_in(reg_psum_23_26), .reg_activation(reg_activation_24_26), .reg_weight(reg_weight_24_26), .reg_partial_sum(reg_psum_24_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_27( .activation_in(reg_activation_24_26), .weight_in(reg_weight_23_27), .partial_sum_in(reg_psum_23_27), .reg_activation(reg_activation_24_27), .reg_weight(reg_weight_24_27), .reg_partial_sum(reg_psum_24_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_28( .activation_in(reg_activation_24_27), .weight_in(reg_weight_23_28), .partial_sum_in(reg_psum_23_28), .reg_activation(reg_activation_24_28), .reg_weight(reg_weight_24_28), .reg_partial_sum(reg_psum_24_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_29( .activation_in(reg_activation_24_28), .weight_in(reg_weight_23_29), .partial_sum_in(reg_psum_23_29), .reg_activation(reg_activation_24_29), .reg_weight(reg_weight_24_29), .reg_partial_sum(reg_psum_24_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_30( .activation_in(reg_activation_24_29), .weight_in(reg_weight_23_30), .partial_sum_in(reg_psum_23_30), .reg_activation(reg_activation_24_30), .reg_weight(reg_weight_24_30), .reg_partial_sum(reg_psum_24_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U24_31( .activation_in(reg_activation_24_30), .weight_in(reg_weight_23_31), .partial_sum_in(reg_psum_23_31), .reg_weight(reg_weight_24_31), .reg_partial_sum(reg_psum_24_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_0( .activation_in(in_activation_25), .weight_in(reg_weight_24_0), .partial_sum_in(reg_psum_24_0), .reg_activation(reg_activation_25_0), .reg_weight(reg_weight_25_0), .reg_partial_sum(reg_psum_25_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_1( .activation_in(reg_activation_25_0), .weight_in(reg_weight_24_1), .partial_sum_in(reg_psum_24_1), .reg_activation(reg_activation_25_1), .reg_weight(reg_weight_25_1), .reg_partial_sum(reg_psum_25_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_2( .activation_in(reg_activation_25_1), .weight_in(reg_weight_24_2), .partial_sum_in(reg_psum_24_2), .reg_activation(reg_activation_25_2), .reg_weight(reg_weight_25_2), .reg_partial_sum(reg_psum_25_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_3( .activation_in(reg_activation_25_2), .weight_in(reg_weight_24_3), .partial_sum_in(reg_psum_24_3), .reg_activation(reg_activation_25_3), .reg_weight(reg_weight_25_3), .reg_partial_sum(reg_psum_25_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_4( .activation_in(reg_activation_25_3), .weight_in(reg_weight_24_4), .partial_sum_in(reg_psum_24_4), .reg_activation(reg_activation_25_4), .reg_weight(reg_weight_25_4), .reg_partial_sum(reg_psum_25_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_5( .activation_in(reg_activation_25_4), .weight_in(reg_weight_24_5), .partial_sum_in(reg_psum_24_5), .reg_activation(reg_activation_25_5), .reg_weight(reg_weight_25_5), .reg_partial_sum(reg_psum_25_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_6( .activation_in(reg_activation_25_5), .weight_in(reg_weight_24_6), .partial_sum_in(reg_psum_24_6), .reg_activation(reg_activation_25_6), .reg_weight(reg_weight_25_6), .reg_partial_sum(reg_psum_25_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_7( .activation_in(reg_activation_25_6), .weight_in(reg_weight_24_7), .partial_sum_in(reg_psum_24_7), .reg_activation(reg_activation_25_7), .reg_weight(reg_weight_25_7), .reg_partial_sum(reg_psum_25_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_8( .activation_in(reg_activation_25_7), .weight_in(reg_weight_24_8), .partial_sum_in(reg_psum_24_8), .reg_activation(reg_activation_25_8), .reg_weight(reg_weight_25_8), .reg_partial_sum(reg_psum_25_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_9( .activation_in(reg_activation_25_8), .weight_in(reg_weight_24_9), .partial_sum_in(reg_psum_24_9), .reg_activation(reg_activation_25_9), .reg_weight(reg_weight_25_9), .reg_partial_sum(reg_psum_25_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_10( .activation_in(reg_activation_25_9), .weight_in(reg_weight_24_10), .partial_sum_in(fault_reg_psum_24_10), .reg_activation(reg_activation_25_10), .reg_weight(reg_weight_25_10), .reg_partial_sum(reg_psum_25_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_11( .activation_in(reg_activation_25_10), .weight_in(reg_weight_24_11), .partial_sum_in(reg_psum_24_11), .reg_activation(reg_activation_25_11), .reg_weight(reg_weight_25_11), .reg_partial_sum(reg_psum_25_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_12( .activation_in(reg_activation_25_11), .weight_in(reg_weight_24_12), .partial_sum_in(reg_psum_24_12), .reg_activation(reg_activation_25_12), .reg_weight(reg_weight_25_12), .reg_partial_sum(reg_psum_25_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_13( .activation_in(reg_activation_25_12), .weight_in(reg_weight_24_13), .partial_sum_in(reg_psum_24_13), .reg_activation(reg_activation_25_13), .reg_weight(reg_weight_25_13), .reg_partial_sum(reg_psum_25_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_14( .activation_in(reg_activation_25_13), .weight_in(reg_weight_24_14), .partial_sum_in(reg_psum_24_14), .reg_activation(reg_activation_25_14), .reg_weight(reg_weight_25_14), .reg_partial_sum(reg_psum_25_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_15( .activation_in(reg_activation_25_14), .weight_in(reg_weight_24_15), .partial_sum_in(reg_psum_24_15), .reg_activation(reg_activation_25_15), .reg_weight(reg_weight_25_15), .reg_partial_sum(reg_psum_25_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_16( .activation_in(reg_activation_25_15), .weight_in(reg_weight_24_16), .partial_sum_in(reg_psum_24_16), .reg_activation(reg_activation_25_16), .reg_weight(reg_weight_25_16), .reg_partial_sum(reg_psum_25_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_17( .activation_in(reg_activation_25_16), .weight_in(reg_weight_24_17), .partial_sum_in(reg_psum_24_17), .reg_activation(reg_activation_25_17), .reg_weight(reg_weight_25_17), .reg_partial_sum(reg_psum_25_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_18( .activation_in(reg_activation_25_17), .weight_in(reg_weight_24_18), .partial_sum_in(reg_psum_24_18), .reg_activation(reg_activation_25_18), .reg_weight(reg_weight_25_18), .reg_partial_sum(reg_psum_25_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_19( .activation_in(reg_activation_25_18), .weight_in(reg_weight_24_19), .partial_sum_in(reg_psum_24_19), .reg_activation(reg_activation_25_19), .reg_weight(reg_weight_25_19), .reg_partial_sum(reg_psum_25_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_20( .activation_in(reg_activation_25_19), .weight_in(reg_weight_24_20), .partial_sum_in(reg_psum_24_20), .reg_activation(reg_activation_25_20), .reg_weight(reg_weight_25_20), .reg_partial_sum(reg_psum_25_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_21( .activation_in(reg_activation_25_20), .weight_in(reg_weight_24_21), .partial_sum_in(reg_psum_24_21), .reg_activation(reg_activation_25_21), .reg_weight(reg_weight_25_21), .reg_partial_sum(reg_psum_25_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_22( .activation_in(reg_activation_25_21), .weight_in(reg_weight_24_22), .partial_sum_in(reg_psum_24_22), .reg_activation(reg_activation_25_22), .reg_weight(reg_weight_25_22), .reg_partial_sum(reg_psum_25_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_23( .activation_in(reg_activation_25_22), .weight_in(reg_weight_24_23), .partial_sum_in(reg_psum_24_23), .reg_activation(reg_activation_25_23), .reg_weight(reg_weight_25_23), .reg_partial_sum(reg_psum_25_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_24( .activation_in(reg_activation_25_23), .weight_in(reg_weight_24_24), .partial_sum_in(reg_psum_24_24), .reg_activation(reg_activation_25_24), .reg_weight(reg_weight_25_24), .reg_partial_sum(reg_psum_25_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_25( .activation_in(reg_activation_25_24), .weight_in(reg_weight_24_25), .partial_sum_in(reg_psum_24_25), .reg_activation(reg_activation_25_25), .reg_weight(reg_weight_25_25), .reg_partial_sum(reg_psum_25_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_26( .activation_in(reg_activation_25_25), .weight_in(reg_weight_24_26), .partial_sum_in(reg_psum_24_26), .reg_activation(reg_activation_25_26), .reg_weight(reg_weight_25_26), .reg_partial_sum(reg_psum_25_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_27( .activation_in(reg_activation_25_26), .weight_in(reg_weight_24_27), .partial_sum_in(reg_psum_24_27), .reg_activation(reg_activation_25_27), .reg_weight(reg_weight_25_27), .reg_partial_sum(reg_psum_25_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_28( .activation_in(reg_activation_25_27), .weight_in(reg_weight_24_28), .partial_sum_in(reg_psum_24_28), .reg_activation(reg_activation_25_28), .reg_weight(reg_weight_25_28), .reg_partial_sum(reg_psum_25_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_29( .activation_in(reg_activation_25_28), .weight_in(reg_weight_24_29), .partial_sum_in(reg_psum_24_29), .reg_activation(reg_activation_25_29), .reg_weight(reg_weight_25_29), .reg_partial_sum(reg_psum_25_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_30( .activation_in(reg_activation_25_29), .weight_in(reg_weight_24_30), .partial_sum_in(reg_psum_24_30), .reg_activation(reg_activation_25_30), .reg_weight(reg_weight_25_30), .reg_partial_sum(reg_psum_25_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U25_31( .activation_in(reg_activation_25_30), .weight_in(reg_weight_24_31), .partial_sum_in(reg_psum_24_31), .reg_weight(reg_weight_25_31), .reg_partial_sum(reg_psum_25_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_0( .activation_in(in_activation_26), .weight_in(reg_weight_25_0), .partial_sum_in(reg_psum_25_0), .reg_activation(reg_activation_26_0), .reg_weight(reg_weight_26_0), .reg_partial_sum(reg_psum_26_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_1( .activation_in(reg_activation_26_0), .weight_in(reg_weight_25_1), .partial_sum_in(reg_psum_25_1), .reg_activation(reg_activation_26_1), .reg_weight(reg_weight_26_1), .reg_partial_sum(reg_psum_26_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_2( .activation_in(reg_activation_26_1), .weight_in(reg_weight_25_2), .partial_sum_in(reg_psum_25_2), .reg_activation(reg_activation_26_2), .reg_weight(reg_weight_26_2), .reg_partial_sum(reg_psum_26_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_3( .activation_in(reg_activation_26_2), .weight_in(reg_weight_25_3), .partial_sum_in(reg_psum_25_3), .reg_activation(reg_activation_26_3), .reg_weight(reg_weight_26_3), .reg_partial_sum(reg_psum_26_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_4( .activation_in(reg_activation_26_3), .weight_in(reg_weight_25_4), .partial_sum_in(reg_psum_25_4), .reg_activation(reg_activation_26_4), .reg_weight(reg_weight_26_4), .reg_partial_sum(reg_psum_26_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_5( .activation_in(reg_activation_26_4), .weight_in(reg_weight_25_5), .partial_sum_in(reg_psum_25_5), .reg_activation(reg_activation_26_5), .reg_weight(reg_weight_26_5), .reg_partial_sum(reg_psum_26_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_6( .activation_in(reg_activation_26_5), .weight_in(reg_weight_25_6), .partial_sum_in(reg_psum_25_6), .reg_activation(reg_activation_26_6), .reg_weight(reg_weight_26_6), .reg_partial_sum(reg_psum_26_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_7( .activation_in(reg_activation_26_6), .weight_in(reg_weight_25_7), .partial_sum_in(reg_psum_25_7), .reg_activation(reg_activation_26_7), .reg_weight(reg_weight_26_7), .reg_partial_sum(reg_psum_26_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_8( .activation_in(reg_activation_26_7), .weight_in(reg_weight_25_8), .partial_sum_in(reg_psum_25_8), .reg_activation(reg_activation_26_8), .reg_weight(reg_weight_26_8), .reg_partial_sum(reg_psum_26_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_9( .activation_in(reg_activation_26_8), .weight_in(reg_weight_25_9), .partial_sum_in(reg_psum_25_9), .reg_activation(reg_activation_26_9), .reg_weight(reg_weight_26_9), .reg_partial_sum(reg_psum_26_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_10( .activation_in(reg_activation_26_9), .weight_in(reg_weight_25_10), .partial_sum_in(reg_psum_25_10), .reg_activation(reg_activation_26_10), .reg_weight(reg_weight_26_10), .reg_partial_sum(reg_psum_26_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_11( .activation_in(reg_activation_26_10), .weight_in(reg_weight_25_11), .partial_sum_in(reg_psum_25_11), .reg_activation(reg_activation_26_11), .reg_weight(reg_weight_26_11), .reg_partial_sum(reg_psum_26_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_12( .activation_in(reg_activation_26_11), .weight_in(reg_weight_25_12), .partial_sum_in(reg_psum_25_12), .reg_activation(reg_activation_26_12), .reg_weight(reg_weight_26_12), .reg_partial_sum(reg_psum_26_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_13( .activation_in(reg_activation_26_12), .weight_in(reg_weight_25_13), .partial_sum_in(reg_psum_25_13), .reg_activation(reg_activation_26_13), .reg_weight(reg_weight_26_13), .reg_partial_sum(reg_psum_26_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_14( .activation_in(reg_activation_26_13), .weight_in(reg_weight_25_14), .partial_sum_in(reg_psum_25_14), .reg_activation(reg_activation_26_14), .reg_weight(reg_weight_26_14), .reg_partial_sum(reg_psum_26_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_15( .activation_in(reg_activation_26_14), .weight_in(reg_weight_25_15), .partial_sum_in(reg_psum_25_15), .reg_activation(reg_activation_26_15), .reg_weight(reg_weight_26_15), .reg_partial_sum(reg_psum_26_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_16( .activation_in(reg_activation_26_15), .weight_in(reg_weight_25_16), .partial_sum_in(reg_psum_25_16), .reg_activation(reg_activation_26_16), .reg_weight(reg_weight_26_16), .reg_partial_sum(reg_psum_26_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_17( .activation_in(reg_activation_26_16), .weight_in(reg_weight_25_17), .partial_sum_in(reg_psum_25_17), .reg_activation(reg_activation_26_17), .reg_weight(reg_weight_26_17), .reg_partial_sum(reg_psum_26_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_18( .activation_in(reg_activation_26_17), .weight_in(reg_weight_25_18), .partial_sum_in(reg_psum_25_18), .reg_activation(reg_activation_26_18), .reg_weight(reg_weight_26_18), .reg_partial_sum(reg_psum_26_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_19( .activation_in(reg_activation_26_18), .weight_in(reg_weight_25_19), .partial_sum_in(reg_psum_25_19), .reg_activation(reg_activation_26_19), .reg_weight(reg_weight_26_19), .reg_partial_sum(reg_psum_26_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_20( .activation_in(reg_activation_26_19), .weight_in(reg_weight_25_20), .partial_sum_in(reg_psum_25_20), .reg_activation(reg_activation_26_20), .reg_weight(reg_weight_26_20), .reg_partial_sum(reg_psum_26_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_21( .activation_in(reg_activation_26_20), .weight_in(reg_weight_25_21), .partial_sum_in(reg_psum_25_21), .reg_activation(reg_activation_26_21), .reg_weight(reg_weight_26_21), .reg_partial_sum(reg_psum_26_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_22( .activation_in(reg_activation_26_21), .weight_in(reg_weight_25_22), .partial_sum_in(reg_psum_25_22), .reg_activation(reg_activation_26_22), .reg_weight(reg_weight_26_22), .reg_partial_sum(reg_psum_26_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_23( .activation_in(reg_activation_26_22), .weight_in(reg_weight_25_23), .partial_sum_in(reg_psum_25_23), .reg_activation(reg_activation_26_23), .reg_weight(reg_weight_26_23), .reg_partial_sum(reg_psum_26_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_24( .activation_in(reg_activation_26_23), .weight_in(reg_weight_25_24), .partial_sum_in(reg_psum_25_24), .reg_activation(reg_activation_26_24), .reg_weight(reg_weight_26_24), .reg_partial_sum(reg_psum_26_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_25( .activation_in(reg_activation_26_24), .weight_in(reg_weight_25_25), .partial_sum_in(reg_psum_25_25), .reg_activation(reg_activation_26_25), .reg_weight(reg_weight_26_25), .reg_partial_sum(reg_psum_26_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_26( .activation_in(reg_activation_26_25), .weight_in(reg_weight_25_26), .partial_sum_in(reg_psum_25_26), .reg_activation(reg_activation_26_26), .reg_weight(reg_weight_26_26), .reg_partial_sum(reg_psum_26_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_27( .activation_in(reg_activation_26_26), .weight_in(reg_weight_25_27), .partial_sum_in(reg_psum_25_27), .reg_activation(reg_activation_26_27), .reg_weight(reg_weight_26_27), .reg_partial_sum(reg_psum_26_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_28( .activation_in(reg_activation_26_27), .weight_in(reg_weight_25_28), .partial_sum_in(reg_psum_25_28), .reg_activation(reg_activation_26_28), .reg_weight(reg_weight_26_28), .reg_partial_sum(reg_psum_26_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_29( .activation_in(reg_activation_26_28), .weight_in(reg_weight_25_29), .partial_sum_in(reg_psum_25_29), .reg_activation(reg_activation_26_29), .reg_weight(reg_weight_26_29), .reg_partial_sum(reg_psum_26_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_30( .activation_in(reg_activation_26_29), .weight_in(reg_weight_25_30), .partial_sum_in(reg_psum_25_30), .reg_activation(reg_activation_26_30), .reg_weight(reg_weight_26_30), .reg_partial_sum(reg_psum_26_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U26_31( .activation_in(reg_activation_26_30), .weight_in(reg_weight_25_31), .partial_sum_in(reg_psum_25_31), .reg_weight(reg_weight_26_31), .reg_partial_sum(reg_psum_26_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_0( .activation_in(in_activation_27), .weight_in(reg_weight_26_0), .partial_sum_in(reg_psum_26_0), .reg_activation(reg_activation_27_0), .reg_weight(reg_weight_27_0), .reg_partial_sum(reg_psum_27_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_1( .activation_in(reg_activation_27_0), .weight_in(reg_weight_26_1), .partial_sum_in(reg_psum_26_1), .reg_activation(reg_activation_27_1), .reg_weight(reg_weight_27_1), .reg_partial_sum(reg_psum_27_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_2( .activation_in(reg_activation_27_1), .weight_in(reg_weight_26_2), .partial_sum_in(reg_psum_26_2), .reg_activation(reg_activation_27_2), .reg_weight(reg_weight_27_2), .reg_partial_sum(reg_psum_27_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_3( .activation_in(reg_activation_27_2), .weight_in(reg_weight_26_3), .partial_sum_in(reg_psum_26_3), .reg_activation(reg_activation_27_3), .reg_weight(reg_weight_27_3), .reg_partial_sum(reg_psum_27_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_4( .activation_in(reg_activation_27_3), .weight_in(reg_weight_26_4), .partial_sum_in(reg_psum_26_4), .reg_activation(reg_activation_27_4), .reg_weight(reg_weight_27_4), .reg_partial_sum(reg_psum_27_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_5( .activation_in(reg_activation_27_4), .weight_in(reg_weight_26_5), .partial_sum_in(reg_psum_26_5), .reg_activation(reg_activation_27_5), .reg_weight(reg_weight_27_5), .reg_partial_sum(reg_psum_27_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_6( .activation_in(reg_activation_27_5), .weight_in(reg_weight_26_6), .partial_sum_in(reg_psum_26_6), .reg_activation(reg_activation_27_6), .reg_weight(reg_weight_27_6), .reg_partial_sum(reg_psum_27_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_7( .activation_in(reg_activation_27_6), .weight_in(reg_weight_26_7), .partial_sum_in(reg_psum_26_7), .reg_activation(reg_activation_27_7), .reg_weight(reg_weight_27_7), .reg_partial_sum(reg_psum_27_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_8( .activation_in(reg_activation_27_7), .weight_in(reg_weight_26_8), .partial_sum_in(reg_psum_26_8), .reg_activation(reg_activation_27_8), .reg_weight(reg_weight_27_8), .reg_partial_sum(reg_psum_27_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_9( .activation_in(reg_activation_27_8), .weight_in(reg_weight_26_9), .partial_sum_in(reg_psum_26_9), .reg_activation(reg_activation_27_9), .reg_weight(reg_weight_27_9), .reg_partial_sum(reg_psum_27_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_10( .activation_in(reg_activation_27_9), .weight_in(reg_weight_26_10), .partial_sum_in(reg_psum_26_10), .reg_activation(reg_activation_27_10), .reg_weight(reg_weight_27_10), .reg_partial_sum(reg_psum_27_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_11( .activation_in(reg_activation_27_10), .weight_in(reg_weight_26_11), .partial_sum_in(reg_psum_26_11), .reg_activation(reg_activation_27_11), .reg_weight(reg_weight_27_11), .reg_partial_sum(reg_psum_27_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_12( .activation_in(reg_activation_27_11), .weight_in(reg_weight_26_12), .partial_sum_in(reg_psum_26_12), .reg_activation(reg_activation_27_12), .reg_weight(reg_weight_27_12), .reg_partial_sum(reg_psum_27_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_13( .activation_in(reg_activation_27_12), .weight_in(reg_weight_26_13), .partial_sum_in(reg_psum_26_13), .reg_activation(reg_activation_27_13), .reg_weight(reg_weight_27_13), .reg_partial_sum(reg_psum_27_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_14( .activation_in(reg_activation_27_13), .weight_in(reg_weight_26_14), .partial_sum_in(reg_psum_26_14), .reg_activation(reg_activation_27_14), .reg_weight(reg_weight_27_14), .reg_partial_sum(reg_psum_27_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_15( .activation_in(reg_activation_27_14), .weight_in(reg_weight_26_15), .partial_sum_in(reg_psum_26_15), .reg_activation(reg_activation_27_15), .reg_weight(reg_weight_27_15), .reg_partial_sum(reg_psum_27_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_16( .activation_in(reg_activation_27_15), .weight_in(reg_weight_26_16), .partial_sum_in(reg_psum_26_16), .reg_activation(reg_activation_27_16), .reg_weight(reg_weight_27_16), .reg_partial_sum(reg_psum_27_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_17( .activation_in(reg_activation_27_16), .weight_in(reg_weight_26_17), .partial_sum_in(reg_psum_26_17), .reg_activation(reg_activation_27_17), .reg_weight(reg_weight_27_17), .reg_partial_sum(reg_psum_27_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_18( .activation_in(reg_activation_27_17), .weight_in(reg_weight_26_18), .partial_sum_in(reg_psum_26_18), .reg_activation(reg_activation_27_18), .reg_weight(reg_weight_27_18), .reg_partial_sum(reg_psum_27_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_19( .activation_in(reg_activation_27_18), .weight_in(reg_weight_26_19), .partial_sum_in(reg_psum_26_19), .reg_activation(reg_activation_27_19), .reg_weight(reg_weight_27_19), .reg_partial_sum(reg_psum_27_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_20( .activation_in(reg_activation_27_19), .weight_in(reg_weight_26_20), .partial_sum_in(reg_psum_26_20), .reg_activation(reg_activation_27_20), .reg_weight(reg_weight_27_20), .reg_partial_sum(reg_psum_27_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_21( .activation_in(reg_activation_27_20), .weight_in(reg_weight_26_21), .partial_sum_in(reg_psum_26_21), .reg_activation(reg_activation_27_21), .reg_weight(reg_weight_27_21), .reg_partial_sum(reg_psum_27_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_22( .activation_in(reg_activation_27_21), .weight_in(reg_weight_26_22), .partial_sum_in(reg_psum_26_22), .reg_activation(reg_activation_27_22), .reg_weight(reg_weight_27_22), .reg_partial_sum(reg_psum_27_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_23( .activation_in(reg_activation_27_22), .weight_in(reg_weight_26_23), .partial_sum_in(reg_psum_26_23), .reg_activation(reg_activation_27_23), .reg_weight(reg_weight_27_23), .reg_partial_sum(reg_psum_27_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_24( .activation_in(reg_activation_27_23), .weight_in(reg_weight_26_24), .partial_sum_in(reg_psum_26_24), .reg_activation(reg_activation_27_24), .reg_weight(reg_weight_27_24), .reg_partial_sum(reg_psum_27_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_25( .activation_in(reg_activation_27_24), .weight_in(reg_weight_26_25), .partial_sum_in(reg_psum_26_25), .reg_activation(reg_activation_27_25), .reg_weight(reg_weight_27_25), .reg_partial_sum(reg_psum_27_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_26( .activation_in(reg_activation_27_25), .weight_in(reg_weight_26_26), .partial_sum_in(reg_psum_26_26), .reg_activation(reg_activation_27_26), .reg_weight(reg_weight_27_26), .reg_partial_sum(reg_psum_27_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_27( .activation_in(reg_activation_27_26), .weight_in(reg_weight_26_27), .partial_sum_in(reg_psum_26_27), .reg_activation(reg_activation_27_27), .reg_weight(reg_weight_27_27), .reg_partial_sum(reg_psum_27_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_28( .activation_in(reg_activation_27_27), .weight_in(reg_weight_26_28), .partial_sum_in(reg_psum_26_28), .reg_activation(reg_activation_27_28), .reg_weight(reg_weight_27_28), .reg_partial_sum(reg_psum_27_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_29( .activation_in(reg_activation_27_28), .weight_in(reg_weight_26_29), .partial_sum_in(reg_psum_26_29), .reg_activation(reg_activation_27_29), .reg_weight(reg_weight_27_29), .reg_partial_sum(reg_psum_27_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_30( .activation_in(reg_activation_27_29), .weight_in(reg_weight_26_30), .partial_sum_in(reg_psum_26_30), .reg_activation(reg_activation_27_30), .reg_weight(reg_weight_27_30), .reg_partial_sum(reg_psum_27_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U27_31( .activation_in(reg_activation_27_30), .weight_in(reg_weight_26_31), .partial_sum_in(reg_psum_26_31), .reg_weight(reg_weight_27_31), .reg_partial_sum(reg_psum_27_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_0( .activation_in(in_activation_28), .weight_in(reg_weight_27_0), .partial_sum_in(reg_psum_27_0), .reg_activation(reg_activation_28_0), .reg_weight(reg_weight_28_0), .reg_partial_sum(reg_psum_28_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_1( .activation_in(reg_activation_28_0), .weight_in(reg_weight_27_1), .partial_sum_in(reg_psum_27_1), .reg_activation(reg_activation_28_1), .reg_weight(reg_weight_28_1), .reg_partial_sum(reg_psum_28_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_2( .activation_in(reg_activation_28_1), .weight_in(reg_weight_27_2), .partial_sum_in(reg_psum_27_2), .reg_activation(reg_activation_28_2), .reg_weight(reg_weight_28_2), .reg_partial_sum(reg_psum_28_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_3( .activation_in(reg_activation_28_2), .weight_in(reg_weight_27_3), .partial_sum_in(reg_psum_27_3), .reg_activation(reg_activation_28_3), .reg_weight(reg_weight_28_3), .reg_partial_sum(reg_psum_28_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_4( .activation_in(reg_activation_28_3), .weight_in(reg_weight_27_4), .partial_sum_in(reg_psum_27_4), .reg_activation(reg_activation_28_4), .reg_weight(reg_weight_28_4), .reg_partial_sum(reg_psum_28_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_5( .activation_in(reg_activation_28_4), .weight_in(reg_weight_27_5), .partial_sum_in(reg_psum_27_5), .reg_activation(reg_activation_28_5), .reg_weight(reg_weight_28_5), .reg_partial_sum(reg_psum_28_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_6( .activation_in(reg_activation_28_5), .weight_in(reg_weight_27_6), .partial_sum_in(reg_psum_27_6), .reg_activation(reg_activation_28_6), .reg_weight(reg_weight_28_6), .reg_partial_sum(reg_psum_28_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_7( .activation_in(reg_activation_28_6), .weight_in(reg_weight_27_7), .partial_sum_in(reg_psum_27_7), .reg_activation(reg_activation_28_7), .reg_weight(reg_weight_28_7), .reg_partial_sum(reg_psum_28_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_8( .activation_in(reg_activation_28_7), .weight_in(reg_weight_27_8), .partial_sum_in(reg_psum_27_8), .reg_activation(reg_activation_28_8), .reg_weight(reg_weight_28_8), .reg_partial_sum(reg_psum_28_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_9( .activation_in(reg_activation_28_8), .weight_in(reg_weight_27_9), .partial_sum_in(reg_psum_27_9), .reg_activation(reg_activation_28_9), .reg_weight(reg_weight_28_9), .reg_partial_sum(reg_psum_28_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_10( .activation_in(reg_activation_28_9), .weight_in(reg_weight_27_10), .partial_sum_in(reg_psum_27_10), .reg_activation(reg_activation_28_10), .reg_weight(reg_weight_28_10), .reg_partial_sum(reg_psum_28_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_11( .activation_in(reg_activation_28_10), .weight_in(reg_weight_27_11), .partial_sum_in(reg_psum_27_11), .reg_activation(reg_activation_28_11), .reg_weight(reg_weight_28_11), .reg_partial_sum(reg_psum_28_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_12( .activation_in(reg_activation_28_11), .weight_in(reg_weight_27_12), .partial_sum_in(reg_psum_27_12), .reg_activation(reg_activation_28_12), .reg_weight(reg_weight_28_12), .reg_partial_sum(reg_psum_28_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_13( .activation_in(reg_activation_28_12), .weight_in(reg_weight_27_13), .partial_sum_in(reg_psum_27_13), .reg_activation(reg_activation_28_13), .reg_weight(reg_weight_28_13), .reg_partial_sum(reg_psum_28_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_14( .activation_in(reg_activation_28_13), .weight_in(reg_weight_27_14), .partial_sum_in(reg_psum_27_14), .reg_activation(reg_activation_28_14), .reg_weight(reg_weight_28_14), .reg_partial_sum(reg_psum_28_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_15( .activation_in(reg_activation_28_14), .weight_in(reg_weight_27_15), .partial_sum_in(reg_psum_27_15), .reg_activation(reg_activation_28_15), .reg_weight(reg_weight_28_15), .reg_partial_sum(reg_psum_28_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_16( .activation_in(reg_activation_28_15), .weight_in(reg_weight_27_16), .partial_sum_in(reg_psum_27_16), .reg_activation(reg_activation_28_16), .reg_weight(reg_weight_28_16), .reg_partial_sum(reg_psum_28_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_17( .activation_in(reg_activation_28_16), .weight_in(reg_weight_27_17), .partial_sum_in(reg_psum_27_17), .reg_activation(reg_activation_28_17), .reg_weight(reg_weight_28_17), .reg_partial_sum(reg_psum_28_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_18( .activation_in(reg_activation_28_17), .weight_in(reg_weight_27_18), .partial_sum_in(reg_psum_27_18), .reg_activation(reg_activation_28_18), .reg_weight(reg_weight_28_18), .reg_partial_sum(reg_psum_28_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_19( .activation_in(reg_activation_28_18), .weight_in(reg_weight_27_19), .partial_sum_in(reg_psum_27_19), .reg_activation(reg_activation_28_19), .reg_weight(reg_weight_28_19), .reg_partial_sum(reg_psum_28_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_20( .activation_in(reg_activation_28_19), .weight_in(reg_weight_27_20), .partial_sum_in(reg_psum_27_20), .reg_activation(reg_activation_28_20), .reg_weight(reg_weight_28_20), .reg_partial_sum(reg_psum_28_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_21( .activation_in(reg_activation_28_20), .weight_in(reg_weight_27_21), .partial_sum_in(reg_psum_27_21), .reg_activation(reg_activation_28_21), .reg_weight(reg_weight_28_21), .reg_partial_sum(reg_psum_28_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_22( .activation_in(reg_activation_28_21), .weight_in(reg_weight_27_22), .partial_sum_in(reg_psum_27_22), .reg_activation(reg_activation_28_22), .reg_weight(reg_weight_28_22), .reg_partial_sum(reg_psum_28_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_23( .activation_in(reg_activation_28_22), .weight_in(reg_weight_27_23), .partial_sum_in(reg_psum_27_23), .reg_activation(reg_activation_28_23), .reg_weight(reg_weight_28_23), .reg_partial_sum(reg_psum_28_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_24( .activation_in(reg_activation_28_23), .weight_in(reg_weight_27_24), .partial_sum_in(reg_psum_27_24), .reg_activation(reg_activation_28_24), .reg_weight(reg_weight_28_24), .reg_partial_sum(reg_psum_28_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_25( .activation_in(reg_activation_28_24), .weight_in(reg_weight_27_25), .partial_sum_in(reg_psum_27_25), .reg_activation(reg_activation_28_25), .reg_weight(reg_weight_28_25), .reg_partial_sum(reg_psum_28_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_26( .activation_in(reg_activation_28_25), .weight_in(reg_weight_27_26), .partial_sum_in(reg_psum_27_26), .reg_activation(reg_activation_28_26), .reg_weight(reg_weight_28_26), .reg_partial_sum(reg_psum_28_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_27( .activation_in(reg_activation_28_26), .weight_in(reg_weight_27_27), .partial_sum_in(reg_psum_27_27), .reg_activation(reg_activation_28_27), .reg_weight(reg_weight_28_27), .reg_partial_sum(reg_psum_28_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_28( .activation_in(reg_activation_28_27), .weight_in(reg_weight_27_28), .partial_sum_in(reg_psum_27_28), .reg_activation(reg_activation_28_28), .reg_weight(reg_weight_28_28), .reg_partial_sum(reg_psum_28_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_29( .activation_in(reg_activation_28_28), .weight_in(reg_weight_27_29), .partial_sum_in(reg_psum_27_29), .reg_activation(reg_activation_28_29), .reg_weight(reg_weight_28_29), .reg_partial_sum(reg_psum_28_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_30( .activation_in(reg_activation_28_29), .weight_in(reg_weight_27_30), .partial_sum_in(reg_psum_27_30), .reg_activation(reg_activation_28_30), .reg_weight(reg_weight_28_30), .reg_partial_sum(reg_psum_28_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U28_31( .activation_in(reg_activation_28_30), .weight_in(reg_weight_27_31), .partial_sum_in(reg_psum_27_31), .reg_weight(reg_weight_28_31), .reg_partial_sum(reg_psum_28_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_0( .activation_in(in_activation_29), .weight_in(reg_weight_28_0), .partial_sum_in(reg_psum_28_0), .reg_activation(reg_activation_29_0), .reg_weight(reg_weight_29_0), .reg_partial_sum(reg_psum_29_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_1( .activation_in(reg_activation_29_0), .weight_in(reg_weight_28_1), .partial_sum_in(reg_psum_28_1), .reg_activation(reg_activation_29_1), .reg_weight(reg_weight_29_1), .reg_partial_sum(reg_psum_29_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_2( .activation_in(reg_activation_29_1), .weight_in(reg_weight_28_2), .partial_sum_in(reg_psum_28_2), .reg_activation(reg_activation_29_2), .reg_weight(reg_weight_29_2), .reg_partial_sum(reg_psum_29_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_3( .activation_in(reg_activation_29_2), .weight_in(reg_weight_28_3), .partial_sum_in(reg_psum_28_3), .reg_activation(reg_activation_29_3), .reg_weight(reg_weight_29_3), .reg_partial_sum(reg_psum_29_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_4( .activation_in(reg_activation_29_3), .weight_in(reg_weight_28_4), .partial_sum_in(reg_psum_28_4), .reg_activation(reg_activation_29_4), .reg_weight(reg_weight_29_4), .reg_partial_sum(reg_psum_29_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_5( .activation_in(reg_activation_29_4), .weight_in(reg_weight_28_5), .partial_sum_in(reg_psum_28_5), .reg_activation(reg_activation_29_5), .reg_weight(reg_weight_29_5), .reg_partial_sum(reg_psum_29_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_6( .activation_in(reg_activation_29_5), .weight_in(reg_weight_28_6), .partial_sum_in(reg_psum_28_6), .reg_activation(reg_activation_29_6), .reg_weight(reg_weight_29_6), .reg_partial_sum(reg_psum_29_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_7( .activation_in(reg_activation_29_6), .weight_in(reg_weight_28_7), .partial_sum_in(reg_psum_28_7), .reg_activation(reg_activation_29_7), .reg_weight(reg_weight_29_7), .reg_partial_sum(reg_psum_29_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_8( .activation_in(reg_activation_29_7), .weight_in(reg_weight_28_8), .partial_sum_in(reg_psum_28_8), .reg_activation(reg_activation_29_8), .reg_weight(reg_weight_29_8), .reg_partial_sum(reg_psum_29_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_9( .activation_in(reg_activation_29_8), .weight_in(reg_weight_28_9), .partial_sum_in(reg_psum_28_9), .reg_activation(reg_activation_29_9), .reg_weight(reg_weight_29_9), .reg_partial_sum(reg_psum_29_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_10( .activation_in(reg_activation_29_9), .weight_in(reg_weight_28_10), .partial_sum_in(reg_psum_28_10), .reg_activation(reg_activation_29_10), .reg_weight(reg_weight_29_10), .reg_partial_sum(reg_psum_29_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_11( .activation_in(reg_activation_29_10), .weight_in(reg_weight_28_11), .partial_sum_in(reg_psum_28_11), .reg_activation(reg_activation_29_11), .reg_weight(reg_weight_29_11), .reg_partial_sum(reg_psum_29_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_12( .activation_in(reg_activation_29_11), .weight_in(reg_weight_28_12), .partial_sum_in(reg_psum_28_12), .reg_activation(reg_activation_29_12), .reg_weight(reg_weight_29_12), .reg_partial_sum(reg_psum_29_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_13( .activation_in(reg_activation_29_12), .weight_in(reg_weight_28_13), .partial_sum_in(reg_psum_28_13), .reg_activation(reg_activation_29_13), .reg_weight(reg_weight_29_13), .reg_partial_sum(reg_psum_29_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_14( .activation_in(reg_activation_29_13), .weight_in(reg_weight_28_14), .partial_sum_in(reg_psum_28_14), .reg_activation(reg_activation_29_14), .reg_weight(reg_weight_29_14), .reg_partial_sum(reg_psum_29_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_15( .activation_in(reg_activation_29_14), .weight_in(reg_weight_28_15), .partial_sum_in(reg_psum_28_15), .reg_activation(reg_activation_29_15), .reg_weight(reg_weight_29_15), .reg_partial_sum(reg_psum_29_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_16( .activation_in(reg_activation_29_15), .weight_in(reg_weight_28_16), .partial_sum_in(reg_psum_28_16), .reg_activation(reg_activation_29_16), .reg_weight(reg_weight_29_16), .reg_partial_sum(reg_psum_29_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_17( .activation_in(reg_activation_29_16), .weight_in(reg_weight_28_17), .partial_sum_in(reg_psum_28_17), .reg_activation(reg_activation_29_17), .reg_weight(reg_weight_29_17), .reg_partial_sum(reg_psum_29_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_18( .activation_in(reg_activation_29_17), .weight_in(reg_weight_28_18), .partial_sum_in(reg_psum_28_18), .reg_activation(reg_activation_29_18), .reg_weight(reg_weight_29_18), .reg_partial_sum(reg_psum_29_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_19( .activation_in(reg_activation_29_18), .weight_in(reg_weight_28_19), .partial_sum_in(reg_psum_28_19), .reg_activation(reg_activation_29_19), .reg_weight(reg_weight_29_19), .reg_partial_sum(reg_psum_29_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_20( .activation_in(reg_activation_29_19), .weight_in(reg_weight_28_20), .partial_sum_in(reg_psum_28_20), .reg_activation(reg_activation_29_20), .reg_weight(reg_weight_29_20), .reg_partial_sum(reg_psum_29_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_21( .activation_in(reg_activation_29_20), .weight_in(reg_weight_28_21), .partial_sum_in(reg_psum_28_21), .reg_activation(reg_activation_29_21), .reg_weight(reg_weight_29_21), .reg_partial_sum(reg_psum_29_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_22( .activation_in(reg_activation_29_21), .weight_in(reg_weight_28_22), .partial_sum_in(reg_psum_28_22), .reg_activation(reg_activation_29_22), .reg_weight(reg_weight_29_22), .reg_partial_sum(reg_psum_29_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_23( .activation_in(reg_activation_29_22), .weight_in(reg_weight_28_23), .partial_sum_in(reg_psum_28_23), .reg_activation(reg_activation_29_23), .reg_weight(reg_weight_29_23), .reg_partial_sum(reg_psum_29_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_24( .activation_in(reg_activation_29_23), .weight_in(reg_weight_28_24), .partial_sum_in(reg_psum_28_24), .reg_activation(reg_activation_29_24), .reg_weight(reg_weight_29_24), .reg_partial_sum(reg_psum_29_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_25( .activation_in(reg_activation_29_24), .weight_in(reg_weight_28_25), .partial_sum_in(reg_psum_28_25), .reg_activation(reg_activation_29_25), .reg_weight(reg_weight_29_25), .reg_partial_sum(reg_psum_29_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_26( .activation_in(reg_activation_29_25), .weight_in(reg_weight_28_26), .partial_sum_in(reg_psum_28_26), .reg_activation(reg_activation_29_26), .reg_weight(reg_weight_29_26), .reg_partial_sum(reg_psum_29_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_27( .activation_in(reg_activation_29_26), .weight_in(reg_weight_28_27), .partial_sum_in(reg_psum_28_27), .reg_activation(reg_activation_29_27), .reg_weight(reg_weight_29_27), .reg_partial_sum(reg_psum_29_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_28( .activation_in(reg_activation_29_27), .weight_in(reg_weight_28_28), .partial_sum_in(reg_psum_28_28), .reg_activation(reg_activation_29_28), .reg_weight(reg_weight_29_28), .reg_partial_sum(reg_psum_29_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_29( .activation_in(reg_activation_29_28), .weight_in(reg_weight_28_29), .partial_sum_in(reg_psum_28_29), .reg_activation(reg_activation_29_29), .reg_weight(reg_weight_29_29), .reg_partial_sum(reg_psum_29_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_30( .activation_in(reg_activation_29_29), .weight_in(reg_weight_28_30), .partial_sum_in(reg_psum_28_30), .reg_activation(reg_activation_29_30), .reg_weight(reg_weight_29_30), .reg_partial_sum(reg_psum_29_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U29_31( .activation_in(reg_activation_29_30), .weight_in(reg_weight_28_31), .partial_sum_in(reg_psum_28_31), .reg_weight(reg_weight_29_31), .reg_partial_sum(reg_psum_29_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_0( .activation_in(in_activation_30), .weight_in(reg_weight_29_0), .partial_sum_in(reg_psum_29_0), .reg_activation(reg_activation_30_0), .reg_weight(reg_weight_30_0), .reg_partial_sum(reg_psum_30_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_1( .activation_in(reg_activation_30_0), .weight_in(reg_weight_29_1), .partial_sum_in(reg_psum_29_1), .reg_activation(reg_activation_30_1), .reg_weight(reg_weight_30_1), .reg_partial_sum(reg_psum_30_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_2( .activation_in(reg_activation_30_1), .weight_in(reg_weight_29_2), .partial_sum_in(reg_psum_29_2), .reg_activation(reg_activation_30_2), .reg_weight(reg_weight_30_2), .reg_partial_sum(reg_psum_30_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_3( .activation_in(reg_activation_30_2), .weight_in(reg_weight_29_3), .partial_sum_in(reg_psum_29_3), .reg_activation(reg_activation_30_3), .reg_weight(reg_weight_30_3), .reg_partial_sum(reg_psum_30_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_4( .activation_in(reg_activation_30_3), .weight_in(reg_weight_29_4), .partial_sum_in(reg_psum_29_4), .reg_activation(reg_activation_30_4), .reg_weight(reg_weight_30_4), .reg_partial_sum(reg_psum_30_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_5( .activation_in(reg_activation_30_4), .weight_in(reg_weight_29_5), .partial_sum_in(reg_psum_29_5), .reg_activation(reg_activation_30_5), .reg_weight(reg_weight_30_5), .reg_partial_sum(reg_psum_30_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_6( .activation_in(reg_activation_30_5), .weight_in(reg_weight_29_6), .partial_sum_in(reg_psum_29_6), .reg_activation(reg_activation_30_6), .reg_weight(reg_weight_30_6), .reg_partial_sum(reg_psum_30_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_7( .activation_in(reg_activation_30_6), .weight_in(reg_weight_29_7), .partial_sum_in(reg_psum_29_7), .reg_activation(reg_activation_30_7), .reg_weight(reg_weight_30_7), .reg_partial_sum(reg_psum_30_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_8( .activation_in(reg_activation_30_7), .weight_in(reg_weight_29_8), .partial_sum_in(reg_psum_29_8), .reg_activation(reg_activation_30_8), .reg_weight(reg_weight_30_8), .reg_partial_sum(reg_psum_30_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_9( .activation_in(reg_activation_30_8), .weight_in(reg_weight_29_9), .partial_sum_in(reg_psum_29_9), .reg_activation(reg_activation_30_9), .reg_weight(reg_weight_30_9), .reg_partial_sum(reg_psum_30_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_10( .activation_in(reg_activation_30_9), .weight_in(reg_weight_29_10), .partial_sum_in(reg_psum_29_10), .reg_activation(reg_activation_30_10), .reg_weight(reg_weight_30_10), .reg_partial_sum(reg_psum_30_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_11( .activation_in(reg_activation_30_10), .weight_in(reg_weight_29_11), .partial_sum_in(reg_psum_29_11), .reg_activation(reg_activation_30_11), .reg_weight(reg_weight_30_11), .reg_partial_sum(reg_psum_30_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_12( .activation_in(reg_activation_30_11), .weight_in(reg_weight_29_12), .partial_sum_in(reg_psum_29_12), .reg_activation(reg_activation_30_12), .reg_weight(reg_weight_30_12), .reg_partial_sum(reg_psum_30_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_13( .activation_in(reg_activation_30_12), .weight_in(reg_weight_29_13), .partial_sum_in(reg_psum_29_13), .reg_activation(reg_activation_30_13), .reg_weight(reg_weight_30_13), .reg_partial_sum(reg_psum_30_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_14( .activation_in(reg_activation_30_13), .weight_in(reg_weight_29_14), .partial_sum_in(reg_psum_29_14), .reg_activation(reg_activation_30_14), .reg_weight(reg_weight_30_14), .reg_partial_sum(reg_psum_30_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_15( .activation_in(reg_activation_30_14), .weight_in(reg_weight_29_15), .partial_sum_in(reg_psum_29_15), .reg_activation(reg_activation_30_15), .reg_weight(reg_weight_30_15), .reg_partial_sum(reg_psum_30_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_16( .activation_in(reg_activation_30_15), .weight_in(reg_weight_29_16), .partial_sum_in(reg_psum_29_16), .reg_activation(reg_activation_30_16), .reg_weight(reg_weight_30_16), .reg_partial_sum(reg_psum_30_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_17( .activation_in(reg_activation_30_16), .weight_in(reg_weight_29_17), .partial_sum_in(reg_psum_29_17), .reg_activation(reg_activation_30_17), .reg_weight(reg_weight_30_17), .reg_partial_sum(reg_psum_30_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_18( .activation_in(reg_activation_30_17), .weight_in(reg_weight_29_18), .partial_sum_in(reg_psum_29_18), .reg_activation(reg_activation_30_18), .reg_weight(reg_weight_30_18), .reg_partial_sum(reg_psum_30_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_19( .activation_in(reg_activation_30_18), .weight_in(reg_weight_29_19), .partial_sum_in(reg_psum_29_19), .reg_activation(reg_activation_30_19), .reg_weight(reg_weight_30_19), .reg_partial_sum(reg_psum_30_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_20( .activation_in(reg_activation_30_19), .weight_in(reg_weight_29_20), .partial_sum_in(reg_psum_29_20), .reg_activation(reg_activation_30_20), .reg_weight(reg_weight_30_20), .reg_partial_sum(reg_psum_30_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_21( .activation_in(reg_activation_30_20), .weight_in(reg_weight_29_21), .partial_sum_in(reg_psum_29_21), .reg_activation(reg_activation_30_21), .reg_weight(reg_weight_30_21), .reg_partial_sum(reg_psum_30_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_22( .activation_in(reg_activation_30_21), .weight_in(reg_weight_29_22), .partial_sum_in(reg_psum_29_22), .reg_activation(reg_activation_30_22), .reg_weight(reg_weight_30_22), .reg_partial_sum(reg_psum_30_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_23( .activation_in(reg_activation_30_22), .weight_in(reg_weight_29_23), .partial_sum_in(reg_psum_29_23), .reg_activation(reg_activation_30_23), .reg_weight(reg_weight_30_23), .reg_partial_sum(reg_psum_30_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_24( .activation_in(reg_activation_30_23), .weight_in(reg_weight_29_24), .partial_sum_in(reg_psum_29_24), .reg_activation(reg_activation_30_24), .reg_weight(reg_weight_30_24), .reg_partial_sum(reg_psum_30_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_25( .activation_in(reg_activation_30_24), .weight_in(reg_weight_29_25), .partial_sum_in(reg_psum_29_25), .reg_activation(reg_activation_30_25), .reg_weight(reg_weight_30_25), .reg_partial_sum(reg_psum_30_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_26( .activation_in(reg_activation_30_25), .weight_in(reg_weight_29_26), .partial_sum_in(reg_psum_29_26), .reg_activation(reg_activation_30_26), .reg_weight(reg_weight_30_26), .reg_partial_sum(reg_psum_30_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_27( .activation_in(reg_activation_30_26), .weight_in(reg_weight_29_27), .partial_sum_in(reg_psum_29_27), .reg_activation(reg_activation_30_27), .reg_weight(reg_weight_30_27), .reg_partial_sum(reg_psum_30_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_28( .activation_in(reg_activation_30_27), .weight_in(reg_weight_29_28), .partial_sum_in(reg_psum_29_28), .reg_activation(reg_activation_30_28), .reg_weight(reg_weight_30_28), .reg_partial_sum(reg_psum_30_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_29( .activation_in(reg_activation_30_28), .weight_in(reg_weight_29_29), .partial_sum_in(reg_psum_29_29), .reg_activation(reg_activation_30_29), .reg_weight(reg_weight_30_29), .reg_partial_sum(reg_psum_30_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_30( .activation_in(reg_activation_30_29), .weight_in(reg_weight_29_30), .partial_sum_in(reg_psum_29_30), .reg_activation(reg_activation_30_30), .reg_weight(reg_weight_30_30), .reg_partial_sum(reg_psum_30_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U30_31( .activation_in(reg_activation_30_30), .weight_in(reg_weight_29_31), .partial_sum_in(reg_psum_29_31), .reg_weight(reg_weight_30_31), .reg_partial_sum(reg_psum_30_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_0( .activation_in(in_activation_31), .weight_in(reg_weight_30_0), .partial_sum_in(reg_psum_30_0), .reg_activation(reg_activation_31_0), .reg_partial_sum(reg_psum_31_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_1( .activation_in(reg_activation_31_0), .weight_in(reg_weight_30_1), .partial_sum_in(reg_psum_30_1), .reg_activation(reg_activation_31_1), .reg_partial_sum(reg_psum_31_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_2( .activation_in(reg_activation_31_1), .weight_in(reg_weight_30_2), .partial_sum_in(reg_psum_30_2), .reg_activation(reg_activation_31_2), .reg_partial_sum(reg_psum_31_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_3( .activation_in(reg_activation_31_2), .weight_in(reg_weight_30_3), .partial_sum_in(reg_psum_30_3), .reg_activation(reg_activation_31_3), .reg_partial_sum(reg_psum_31_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_4( .activation_in(reg_activation_31_3), .weight_in(reg_weight_30_4), .partial_sum_in(reg_psum_30_4), .reg_activation(reg_activation_31_4), .reg_partial_sum(reg_psum_31_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_5( .activation_in(reg_activation_31_4), .weight_in(reg_weight_30_5), .partial_sum_in(reg_psum_30_5), .reg_activation(reg_activation_31_5), .reg_partial_sum(reg_psum_31_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_6( .activation_in(reg_activation_31_5), .weight_in(reg_weight_30_6), .partial_sum_in(reg_psum_30_6), .reg_activation(reg_activation_31_6), .reg_partial_sum(reg_psum_31_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_7( .activation_in(reg_activation_31_6), .weight_in(reg_weight_30_7), .partial_sum_in(reg_psum_30_7), .reg_activation(reg_activation_31_7), .reg_partial_sum(reg_psum_31_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_8( .activation_in(reg_activation_31_7), .weight_in(reg_weight_30_8), .partial_sum_in(reg_psum_30_8), .reg_activation(reg_activation_31_8), .reg_partial_sum(reg_psum_31_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_9( .activation_in(reg_activation_31_8), .weight_in(reg_weight_30_9), .partial_sum_in(reg_psum_30_9), .reg_activation(reg_activation_31_9), .reg_partial_sum(reg_psum_31_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_10( .activation_in(reg_activation_31_9), .weight_in(reg_weight_30_10), .partial_sum_in(reg_psum_30_10), .reg_activation(reg_activation_31_10), .reg_partial_sum(reg_psum_31_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_11( .activation_in(reg_activation_31_10), .weight_in(reg_weight_30_11), .partial_sum_in(fault_reg_psum_30_11), .reg_activation(reg_activation_31_11), .reg_partial_sum(reg_psum_31_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_12( .activation_in(reg_activation_31_11), .weight_in(reg_weight_30_12), .partial_sum_in(reg_psum_30_12), .reg_activation(reg_activation_31_12), .reg_partial_sum(reg_psum_31_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_13( .activation_in(reg_activation_31_12), .weight_in(reg_weight_30_13), .partial_sum_in(reg_psum_30_13), .reg_activation(reg_activation_31_13), .reg_partial_sum(reg_psum_31_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_14( .activation_in(reg_activation_31_13), .weight_in(reg_weight_30_14), .partial_sum_in(reg_psum_30_14), .reg_activation(reg_activation_31_14), .reg_partial_sum(reg_psum_31_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_15( .activation_in(reg_activation_31_14), .weight_in(reg_weight_30_15), .partial_sum_in(reg_psum_30_15), .reg_activation(reg_activation_31_15), .reg_partial_sum(reg_psum_31_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_16( .activation_in(reg_activation_31_15), .weight_in(reg_weight_30_16), .partial_sum_in(reg_psum_30_16), .reg_activation(reg_activation_31_16), .reg_partial_sum(reg_psum_31_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_17( .activation_in(reg_activation_31_16), .weight_in(reg_weight_30_17), .partial_sum_in(reg_psum_30_17), .reg_activation(reg_activation_31_17), .reg_partial_sum(reg_psum_31_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_18( .activation_in(reg_activation_31_17), .weight_in(reg_weight_30_18), .partial_sum_in(reg_psum_30_18), .reg_activation(reg_activation_31_18), .reg_partial_sum(reg_psum_31_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_19( .activation_in(reg_activation_31_18), .weight_in(reg_weight_30_19), .partial_sum_in(reg_psum_30_19), .reg_activation(reg_activation_31_19), .reg_partial_sum(reg_psum_31_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_20( .activation_in(reg_activation_31_19), .weight_in(reg_weight_30_20), .partial_sum_in(reg_psum_30_20), .reg_activation(reg_activation_31_20), .reg_partial_sum(reg_psum_31_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_21( .activation_in(reg_activation_31_20), .weight_in(reg_weight_30_21), .partial_sum_in(reg_psum_30_21), .reg_activation(reg_activation_31_21), .reg_partial_sum(reg_psum_31_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_22( .activation_in(reg_activation_31_21), .weight_in(reg_weight_30_22), .partial_sum_in(reg_psum_30_22), .reg_activation(reg_activation_31_22), .reg_partial_sum(reg_psum_31_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_23( .activation_in(reg_activation_31_22), .weight_in(reg_weight_30_23), .partial_sum_in(reg_psum_30_23), .reg_activation(reg_activation_31_23), .reg_partial_sum(reg_psum_31_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_24( .activation_in(reg_activation_31_23), .weight_in(reg_weight_30_24), .partial_sum_in(reg_psum_30_24), .reg_activation(reg_activation_31_24), .reg_partial_sum(reg_psum_31_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_25( .activation_in(reg_activation_31_24), .weight_in(reg_weight_30_25), .partial_sum_in(reg_psum_30_25), .reg_activation(reg_activation_31_25), .reg_partial_sum(reg_psum_31_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_26( .activation_in(reg_activation_31_25), .weight_in(reg_weight_30_26), .partial_sum_in(reg_psum_30_26), .reg_activation(reg_activation_31_26), .reg_partial_sum(reg_psum_31_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_27( .activation_in(reg_activation_31_26), .weight_in(reg_weight_30_27), .partial_sum_in(reg_psum_30_27), .reg_activation(reg_activation_31_27), .reg_partial_sum(reg_psum_31_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_28( .activation_in(reg_activation_31_27), .weight_in(reg_weight_30_28), .partial_sum_in(reg_psum_30_28), .reg_activation(reg_activation_31_28), .reg_partial_sum(reg_psum_31_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_29( .activation_in(reg_activation_31_28), .weight_in(reg_weight_30_29), .partial_sum_in(reg_psum_30_29), .reg_activation(reg_activation_31_29), .reg_partial_sum(reg_psum_31_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_30( .activation_in(reg_activation_31_29), .weight_in(reg_weight_30_30), .partial_sum_in(reg_psum_30_30), .reg_activation(reg_activation_31_30), .reg_partial_sum(reg_psum_31_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE U31_31( .activation_in(reg_activation_31_30), .weight_in(reg_weight_30_31), .partial_sum_in(reg_psum_30_31), .reg_partial_sum(reg_psum_31_31), .clk(clk), .rst(rst), .weight_en(weight_en));
wire signed[15:0]    spare_reg_activation_0_0;
wire signed[15:0]    spare_reg_activation_0_1;
wire signed[15:0]    spare_reg_activation_0_2;
wire signed[15:0]    spare_reg_activation_0_3;
wire signed[15:0]    spare_reg_activation_0_4;
wire signed[15:0]    spare_reg_activation_0_5;
wire signed[15:0]    spare_reg_activation_0_6;
wire signed[15:0]    spare_reg_activation_0_7;
wire signed[15:0]    spare_reg_activation_0_8;
wire signed[15:0]    spare_reg_activation_0_9;
wire signed[15:0]    spare_reg_activation_0_10;
wire signed[15:0]    spare_reg_activation_0_11;
wire signed[15:0]    spare_reg_activation_0_12;
wire signed[15:0]    spare_reg_activation_0_13;
wire signed[15:0]    spare_reg_activation_0_14;
wire signed[15:0]    spare_reg_activation_0_15;
wire signed[15:0]    spare_reg_activation_0_16;
wire signed[15:0]    spare_reg_activation_0_17;
wire signed[15:0]    spare_reg_activation_0_18;
wire signed[15:0]    spare_reg_activation_0_19;
wire signed[15:0]    spare_reg_activation_0_20;
wire signed[15:0]    spare_reg_activation_0_21;
wire signed[15:0]    spare_reg_activation_0_22;
wire signed[15:0]    spare_reg_activation_0_23;
wire signed[15:0]    spare_reg_activation_0_24;
wire signed[15:0]    spare_reg_activation_0_25;
wire signed[15:0]    spare_reg_activation_0_26;
wire signed[15:0]    spare_reg_activation_0_27;
wire signed[15:0]    spare_reg_activation_0_28;
wire signed[15:0]    spare_reg_activation_0_29;
wire signed[15:0]    spare_reg_activation_0_30;
wire signed[15:0]    spare_reg_activation_0_31;
wire signed[15:0]    spare_reg_activation_1_0;
wire signed[15:0]    spare_reg_activation_1_1;
wire signed[15:0]    spare_reg_activation_1_2;
wire signed[15:0]    spare_reg_activation_1_3;
wire signed[15:0]    spare_reg_activation_1_4;
wire signed[15:0]    spare_reg_activation_1_5;
wire signed[15:0]    spare_reg_activation_1_6;
wire signed[15:0]    spare_reg_activation_1_7;
wire signed[15:0]    spare_reg_activation_1_8;
wire signed[15:0]    spare_reg_activation_1_9;
wire signed[15:0]    spare_reg_activation_1_10;
wire signed[15:0]    spare_reg_activation_1_11;
wire signed[15:0]    spare_reg_activation_1_12;
wire signed[15:0]    spare_reg_activation_1_13;
wire signed[15:0]    spare_reg_activation_1_14;
wire signed[15:0]    spare_reg_activation_1_15;
wire signed[15:0]    spare_reg_activation_1_16;
wire signed[15:0]    spare_reg_activation_1_17;
wire signed[15:0]    spare_reg_activation_1_18;
wire signed[15:0]    spare_reg_activation_1_19;
wire signed[15:0]    spare_reg_activation_1_20;
wire signed[15:0]    spare_reg_activation_1_21;
wire signed[15:0]    spare_reg_activation_1_22;
wire signed[15:0]    spare_reg_activation_1_23;
wire signed[15:0]    spare_reg_activation_1_24;
wire signed[15:0]    spare_reg_activation_1_25;
wire signed[15:0]    spare_reg_activation_1_26;
wire signed[15:0]    spare_reg_activation_1_27;
wire signed[15:0]    spare_reg_activation_1_28;
wire signed[15:0]    spare_reg_activation_1_29;
wire signed[15:0]    spare_reg_activation_1_30;
wire signed[15:0]    spare_reg_activation_1_31;
wire signed[15:0]    spare_reg_activation_2_0;
wire signed[15:0]    spare_reg_activation_2_1;
wire signed[15:0]    spare_reg_activation_2_2;
wire signed[15:0]    spare_reg_activation_2_3;
wire signed[15:0]    spare_reg_activation_2_4;
wire signed[15:0]    spare_reg_activation_2_5;
wire signed[15:0]    spare_reg_activation_2_6;
wire signed[15:0]    spare_reg_activation_2_7;
wire signed[15:0]    spare_reg_activation_2_8;
wire signed[15:0]    spare_reg_activation_2_9;
wire signed[15:0]    spare_reg_activation_2_10;
wire signed[15:0]    spare_reg_activation_2_11;
wire signed[15:0]    spare_reg_activation_2_12;
wire signed[15:0]    spare_reg_activation_2_13;
wire signed[15:0]    spare_reg_activation_2_14;
wire signed[15:0]    spare_reg_activation_2_15;
wire signed[15:0]    spare_reg_activation_2_16;
wire signed[15:0]    spare_reg_activation_2_17;
wire signed[15:0]    spare_reg_activation_2_18;
wire signed[15:0]    spare_reg_activation_2_19;
wire signed[15:0]    spare_reg_activation_2_20;
wire signed[15:0]    spare_reg_activation_2_21;
wire signed[15:0]    spare_reg_activation_2_22;
wire signed[15:0]    spare_reg_activation_2_23;
wire signed[15:0]    spare_reg_activation_2_24;
wire signed[15:0]    spare_reg_activation_2_25;
wire signed[15:0]    spare_reg_activation_2_26;
wire signed[15:0]    spare_reg_activation_2_27;
wire signed[15:0]    spare_reg_activation_2_28;
wire signed[15:0]    spare_reg_activation_2_29;
wire signed[15:0]    spare_reg_activation_2_30;
wire signed[15:0]    spare_reg_activation_2_31;
wire signed[15:0]    spare_reg_activation_3_0;
wire signed[15:0]    spare_reg_activation_3_1;
wire signed[15:0]    spare_reg_activation_3_2;
wire signed[15:0]    spare_reg_activation_3_3;
wire signed[15:0]    spare_reg_activation_3_4;
wire signed[15:0]    spare_reg_activation_3_5;
wire signed[15:0]    spare_reg_activation_3_6;
wire signed[15:0]    spare_reg_activation_3_7;
wire signed[15:0]    spare_reg_activation_3_8;
wire signed[15:0]    spare_reg_activation_3_9;
wire signed[15:0]    spare_reg_activation_3_10;
wire signed[15:0]    spare_reg_activation_3_11;
wire signed[15:0]    spare_reg_activation_3_12;
wire signed[15:0]    spare_reg_activation_3_13;
wire signed[15:0]    spare_reg_activation_3_14;
wire signed[15:0]    spare_reg_activation_3_15;
wire signed[15:0]    spare_reg_activation_3_16;
wire signed[15:0]    spare_reg_activation_3_17;
wire signed[15:0]    spare_reg_activation_3_18;
wire signed[15:0]    spare_reg_activation_3_19;
wire signed[15:0]    spare_reg_activation_3_20;
wire signed[15:0]    spare_reg_activation_3_21;
wire signed[15:0]    spare_reg_activation_3_22;
wire signed[15:0]    spare_reg_activation_3_23;
wire signed[15:0]    spare_reg_activation_3_24;
wire signed[15:0]    spare_reg_activation_3_25;
wire signed[15:0]    spare_reg_activation_3_26;
wire signed[15:0]    spare_reg_activation_3_27;
wire signed[15:0]    spare_reg_activation_3_28;
wire signed[15:0]    spare_reg_activation_3_29;
wire signed[15:0]    spare_reg_activation_3_30;
wire signed[15:0]    spare_reg_activation_3_31;
wire signed[15:0]    spare_reg_activation_4_0;
wire signed[15:0]    spare_reg_activation_4_1;
wire signed[15:0]    spare_reg_activation_4_2;
wire signed[15:0]    spare_reg_activation_4_3;
wire signed[15:0]    spare_reg_activation_4_4;
wire signed[15:0]    spare_reg_activation_4_5;
wire signed[15:0]    spare_reg_activation_4_6;
wire signed[15:0]    spare_reg_activation_4_7;
wire signed[15:0]    spare_reg_activation_4_8;
wire signed[15:0]    spare_reg_activation_4_9;
wire signed[15:0]    spare_reg_activation_4_10;
wire signed[15:0]    spare_reg_activation_4_11;
wire signed[15:0]    spare_reg_activation_4_12;
wire signed[15:0]    spare_reg_activation_4_13;
wire signed[15:0]    spare_reg_activation_4_14;
wire signed[15:0]    spare_reg_activation_4_15;
wire signed[15:0]    spare_reg_activation_4_16;
wire signed[15:0]    spare_reg_activation_4_17;
wire signed[15:0]    spare_reg_activation_4_18;
wire signed[15:0]    spare_reg_activation_4_19;
wire signed[15:0]    spare_reg_activation_4_20;
wire signed[15:0]    spare_reg_activation_4_21;
wire signed[15:0]    spare_reg_activation_4_22;
wire signed[15:0]    spare_reg_activation_4_23;
wire signed[15:0]    spare_reg_activation_4_24;
wire signed[15:0]    spare_reg_activation_4_25;
wire signed[15:0]    spare_reg_activation_4_26;
wire signed[15:0]    spare_reg_activation_4_27;
wire signed[15:0]    spare_reg_activation_4_28;
wire signed[15:0]    spare_reg_activation_4_29;
wire signed[15:0]    spare_reg_activation_4_30;
wire signed[15:0]    spare_reg_activation_4_31;
wire signed[15:0]    spare_reg_activation_5_0;
wire signed[15:0]    spare_reg_activation_5_1;
wire signed[15:0]    spare_reg_activation_5_2;
wire signed[15:0]    spare_reg_activation_5_3;
wire signed[15:0]    spare_reg_activation_5_4;
wire signed[15:0]    spare_reg_activation_5_5;
wire signed[15:0]    spare_reg_activation_5_6;
wire signed[15:0]    spare_reg_activation_5_7;
wire signed[15:0]    spare_reg_activation_5_8;
wire signed[15:0]    spare_reg_activation_5_9;
wire signed[15:0]    spare_reg_activation_5_10;
wire signed[15:0]    spare_reg_activation_5_11;
wire signed[15:0]    spare_reg_activation_5_12;
wire signed[15:0]    spare_reg_activation_5_13;
wire signed[15:0]    spare_reg_activation_5_14;
wire signed[15:0]    spare_reg_activation_5_15;
wire signed[15:0]    spare_reg_activation_5_16;
wire signed[15:0]    spare_reg_activation_5_17;
wire signed[15:0]    spare_reg_activation_5_18;
wire signed[15:0]    spare_reg_activation_5_19;
wire signed[15:0]    spare_reg_activation_5_20;
wire signed[15:0]    spare_reg_activation_5_21;
wire signed[15:0]    spare_reg_activation_5_22;
wire signed[15:0]    spare_reg_activation_5_23;
wire signed[15:0]    spare_reg_activation_5_24;
wire signed[15:0]    spare_reg_activation_5_25;
wire signed[15:0]    spare_reg_activation_5_26;
wire signed[15:0]    spare_reg_activation_5_27;
wire signed[15:0]    spare_reg_activation_5_28;
wire signed[15:0]    spare_reg_activation_5_29;
wire signed[15:0]    spare_reg_activation_5_30;
wire signed[15:0]    spare_reg_activation_5_31;
wire signed[15:0]    spare_reg_activation_6_0;
wire signed[15:0]    spare_reg_activation_6_1;
wire signed[15:0]    spare_reg_activation_6_2;
wire signed[15:0]    spare_reg_activation_6_3;
wire signed[15:0]    spare_reg_activation_6_4;
wire signed[15:0]    spare_reg_activation_6_5;
wire signed[15:0]    spare_reg_activation_6_6;
wire signed[15:0]    spare_reg_activation_6_7;
wire signed[15:0]    spare_reg_activation_6_8;
wire signed[15:0]    spare_reg_activation_6_9;
wire signed[15:0]    spare_reg_activation_6_10;
wire signed[15:0]    spare_reg_activation_6_11;
wire signed[15:0]    spare_reg_activation_6_12;
wire signed[15:0]    spare_reg_activation_6_13;
wire signed[15:0]    spare_reg_activation_6_14;
wire signed[15:0]    spare_reg_activation_6_15;
wire signed[15:0]    spare_reg_activation_6_16;
wire signed[15:0]    spare_reg_activation_6_17;
wire signed[15:0]    spare_reg_activation_6_18;
wire signed[15:0]    spare_reg_activation_6_19;
wire signed[15:0]    spare_reg_activation_6_20;
wire signed[15:0]    spare_reg_activation_6_21;
wire signed[15:0]    spare_reg_activation_6_22;
wire signed[15:0]    spare_reg_activation_6_23;
wire signed[15:0]    spare_reg_activation_6_24;
wire signed[15:0]    spare_reg_activation_6_25;
wire signed[15:0]    spare_reg_activation_6_26;
wire signed[15:0]    spare_reg_activation_6_27;
wire signed[15:0]    spare_reg_activation_6_28;
wire signed[15:0]    spare_reg_activation_6_29;
wire signed[15:0]    spare_reg_activation_6_30;
wire signed[15:0]    spare_reg_activation_6_31;
wire signed[15:0]    spare_reg_activation_7_0;
wire signed[15:0]    spare_reg_activation_7_1;
wire signed[15:0]    spare_reg_activation_7_2;
wire signed[15:0]    spare_reg_activation_7_3;
wire signed[15:0]    spare_reg_activation_7_4;
wire signed[15:0]    spare_reg_activation_7_5;
wire signed[15:0]    spare_reg_activation_7_6;
wire signed[15:0]    spare_reg_activation_7_7;
wire signed[15:0]    spare_reg_activation_7_8;
wire signed[15:0]    spare_reg_activation_7_9;
wire signed[15:0]    spare_reg_activation_7_10;
wire signed[15:0]    spare_reg_activation_7_11;
wire signed[15:0]    spare_reg_activation_7_12;
wire signed[15:0]    spare_reg_activation_7_13;
wire signed[15:0]    spare_reg_activation_7_14;
wire signed[15:0]    spare_reg_activation_7_15;
wire signed[15:0]    spare_reg_activation_7_16;
wire signed[15:0]    spare_reg_activation_7_17;
wire signed[15:0]    spare_reg_activation_7_18;
wire signed[15:0]    spare_reg_activation_7_19;
wire signed[15:0]    spare_reg_activation_7_20;
wire signed[15:0]    spare_reg_activation_7_21;
wire signed[15:0]    spare_reg_activation_7_22;
wire signed[15:0]    spare_reg_activation_7_23;
wire signed[15:0]    spare_reg_activation_7_24;
wire signed[15:0]    spare_reg_activation_7_25;
wire signed[15:0]    spare_reg_activation_7_26;
wire signed[15:0]    spare_reg_activation_7_27;
wire signed[15:0]    spare_reg_activation_7_28;
wire signed[15:0]    spare_reg_activation_7_29;
wire signed[15:0]    spare_reg_activation_7_30;
wire signed[15:0]    spare_reg_activation_7_31;
wire signed[15:0]    spare_reg_activation_8_0;
wire signed[15:0]    spare_reg_activation_8_1;
wire signed[15:0]    spare_reg_activation_8_2;
wire signed[15:0]    spare_reg_activation_8_3;
wire signed[15:0]    spare_reg_activation_8_4;
wire signed[15:0]    spare_reg_activation_8_5;
wire signed[15:0]    spare_reg_activation_8_6;
wire signed[15:0]    spare_reg_activation_8_7;
wire signed[15:0]    spare_reg_activation_8_8;
wire signed[15:0]    spare_reg_activation_8_9;
wire signed[15:0]    spare_reg_activation_8_10;
wire signed[15:0]    spare_reg_activation_8_11;
wire signed[15:0]    spare_reg_activation_8_12;
wire signed[15:0]    spare_reg_activation_8_13;
wire signed[15:0]    spare_reg_activation_8_14;
wire signed[15:0]    spare_reg_activation_8_15;
wire signed[15:0]    spare_reg_activation_8_16;
wire signed[15:0]    spare_reg_activation_8_17;
wire signed[15:0]    spare_reg_activation_8_18;
wire signed[15:0]    spare_reg_activation_8_19;
wire signed[15:0]    spare_reg_activation_8_20;
wire signed[15:0]    spare_reg_activation_8_21;
wire signed[15:0]    spare_reg_activation_8_22;
wire signed[15:0]    spare_reg_activation_8_23;
wire signed[15:0]    spare_reg_activation_8_24;
wire signed[15:0]    spare_reg_activation_8_25;
wire signed[15:0]    spare_reg_activation_8_26;
wire signed[15:0]    spare_reg_activation_8_27;
wire signed[15:0]    spare_reg_activation_8_28;
wire signed[15:0]    spare_reg_activation_8_29;
wire signed[15:0]    spare_reg_activation_8_30;
wire signed[15:0]    spare_reg_activation_8_31;
wire signed[15:0]    spare_reg_activation_9_0;
wire signed[15:0]    spare_reg_activation_9_1;
wire signed[15:0]    spare_reg_activation_9_2;
wire signed[15:0]    spare_reg_activation_9_3;
wire signed[15:0]    spare_reg_activation_9_4;
wire signed[15:0]    spare_reg_activation_9_5;
wire signed[15:0]    spare_reg_activation_9_6;
wire signed[15:0]    spare_reg_activation_9_7;
wire signed[15:0]    spare_reg_activation_9_8;
wire signed[15:0]    spare_reg_activation_9_9;
wire signed[15:0]    spare_reg_activation_9_10;
wire signed[15:0]    spare_reg_activation_9_11;
wire signed[15:0]    spare_reg_activation_9_12;
wire signed[15:0]    spare_reg_activation_9_13;
wire signed[15:0]    spare_reg_activation_9_14;
wire signed[15:0]    spare_reg_activation_9_15;
wire signed[15:0]    spare_reg_activation_9_16;
wire signed[15:0]    spare_reg_activation_9_17;
wire signed[15:0]    spare_reg_activation_9_18;
wire signed[15:0]    spare_reg_activation_9_19;
wire signed[15:0]    spare_reg_activation_9_20;
wire signed[15:0]    spare_reg_activation_9_21;
wire signed[15:0]    spare_reg_activation_9_22;
wire signed[15:0]    spare_reg_activation_9_23;
wire signed[15:0]    spare_reg_activation_9_24;
wire signed[15:0]    spare_reg_activation_9_25;
wire signed[15:0]    spare_reg_activation_9_26;
wire signed[15:0]    spare_reg_activation_9_27;
wire signed[15:0]    spare_reg_activation_9_28;
wire signed[15:0]    spare_reg_activation_9_29;
wire signed[15:0]    spare_reg_activation_9_30;
wire signed[15:0]    spare_reg_activation_9_31;
wire signed[15:0]    spare_reg_activation_10_0;
wire signed[15:0]    spare_reg_activation_10_1;
wire signed[15:0]    spare_reg_activation_10_2;
wire signed[15:0]    spare_reg_activation_10_3;
wire signed[15:0]    spare_reg_activation_10_4;
wire signed[15:0]    spare_reg_activation_10_5;
wire signed[15:0]    spare_reg_activation_10_6;
wire signed[15:0]    spare_reg_activation_10_7;
wire signed[15:0]    spare_reg_activation_10_8;
wire signed[15:0]    spare_reg_activation_10_9;
wire signed[15:0]    spare_reg_activation_10_10;
wire signed[15:0]    spare_reg_activation_10_11;
wire signed[15:0]    spare_reg_activation_10_12;
wire signed[15:0]    spare_reg_activation_10_13;
wire signed[15:0]    spare_reg_activation_10_14;
wire signed[15:0]    spare_reg_activation_10_15;
wire signed[15:0]    spare_reg_activation_10_16;
wire signed[15:0]    spare_reg_activation_10_17;
wire signed[15:0]    spare_reg_activation_10_18;
wire signed[15:0]    spare_reg_activation_10_19;
wire signed[15:0]    spare_reg_activation_10_20;
wire signed[15:0]    spare_reg_activation_10_21;
wire signed[15:0]    spare_reg_activation_10_22;
wire signed[15:0]    spare_reg_activation_10_23;
wire signed[15:0]    spare_reg_activation_10_24;
wire signed[15:0]    spare_reg_activation_10_25;
wire signed[15:0]    spare_reg_activation_10_26;
wire signed[15:0]    spare_reg_activation_10_27;
wire signed[15:0]    spare_reg_activation_10_28;
wire signed[15:0]    spare_reg_activation_10_29;
wire signed[15:0]    spare_reg_activation_10_30;
wire signed[15:0]    spare_reg_activation_10_31;
wire signed[15:0]    spare_reg_activation_11_0;
wire signed[15:0]    spare_reg_activation_11_1;
wire signed[15:0]    spare_reg_activation_11_2;
wire signed[15:0]    spare_reg_activation_11_3;
wire signed[15:0]    spare_reg_activation_11_4;
wire signed[15:0]    spare_reg_activation_11_5;
wire signed[15:0]    spare_reg_activation_11_6;
wire signed[15:0]    spare_reg_activation_11_7;
wire signed[15:0]    spare_reg_activation_11_8;
wire signed[15:0]    spare_reg_activation_11_9;
wire signed[15:0]    spare_reg_activation_11_10;
wire signed[15:0]    spare_reg_activation_11_11;
wire signed[15:0]    spare_reg_activation_11_12;
wire signed[15:0]    spare_reg_activation_11_13;
wire signed[15:0]    spare_reg_activation_11_14;
wire signed[15:0]    spare_reg_activation_11_15;
wire signed[15:0]    spare_reg_activation_11_16;
wire signed[15:0]    spare_reg_activation_11_17;
wire signed[15:0]    spare_reg_activation_11_18;
wire signed[15:0]    spare_reg_activation_11_19;
wire signed[15:0]    spare_reg_activation_11_20;
wire signed[15:0]    spare_reg_activation_11_21;
wire signed[15:0]    spare_reg_activation_11_22;
wire signed[15:0]    spare_reg_activation_11_23;
wire signed[15:0]    spare_reg_activation_11_24;
wire signed[15:0]    spare_reg_activation_11_25;
wire signed[15:0]    spare_reg_activation_11_26;
wire signed[15:0]    spare_reg_activation_11_27;
wire signed[15:0]    spare_reg_activation_11_28;
wire signed[15:0]    spare_reg_activation_11_29;
wire signed[15:0]    spare_reg_activation_11_30;
wire signed[15:0]    spare_reg_activation_11_31;
wire signed[15:0]    spare_reg_activation_12_0;
wire signed[15:0]    spare_reg_activation_12_1;
wire signed[15:0]    spare_reg_activation_12_2;
wire signed[15:0]    spare_reg_activation_12_3;
wire signed[15:0]    spare_reg_activation_12_4;
wire signed[15:0]    spare_reg_activation_12_5;
wire signed[15:0]    spare_reg_activation_12_6;
wire signed[15:0]    spare_reg_activation_12_7;
wire signed[15:0]    spare_reg_activation_12_8;
wire signed[15:0]    spare_reg_activation_12_9;
wire signed[15:0]    spare_reg_activation_12_10;
wire signed[15:0]    spare_reg_activation_12_11;
wire signed[15:0]    spare_reg_activation_12_12;
wire signed[15:0]    spare_reg_activation_12_13;
wire signed[15:0]    spare_reg_activation_12_14;
wire signed[15:0]    spare_reg_activation_12_15;
wire signed[15:0]    spare_reg_activation_12_16;
wire signed[15:0]    spare_reg_activation_12_17;
wire signed[15:0]    spare_reg_activation_12_18;
wire signed[15:0]    spare_reg_activation_12_19;
wire signed[15:0]    spare_reg_activation_12_20;
wire signed[15:0]    spare_reg_activation_12_21;
wire signed[15:0]    spare_reg_activation_12_22;
wire signed[15:0]    spare_reg_activation_12_23;
wire signed[15:0]    spare_reg_activation_12_24;
wire signed[15:0]    spare_reg_activation_12_25;
wire signed[15:0]    spare_reg_activation_12_26;
wire signed[15:0]    spare_reg_activation_12_27;
wire signed[15:0]    spare_reg_activation_12_28;
wire signed[15:0]    spare_reg_activation_12_29;
wire signed[15:0]    spare_reg_activation_12_30;
wire signed[15:0]    spare_reg_activation_12_31;
wire signed[15:0]    spare_reg_activation_13_0;
wire signed[15:0]    spare_reg_activation_13_1;
wire signed[15:0]    spare_reg_activation_13_2;
wire signed[15:0]    spare_reg_activation_13_3;
wire signed[15:0]    spare_reg_activation_13_4;
wire signed[15:0]    spare_reg_activation_13_5;
wire signed[15:0]    spare_reg_activation_13_6;
wire signed[15:0]    spare_reg_activation_13_7;
wire signed[15:0]    spare_reg_activation_13_8;
wire signed[15:0]    spare_reg_activation_13_9;
wire signed[15:0]    spare_reg_activation_13_10;
wire signed[15:0]    spare_reg_activation_13_11;
wire signed[15:0]    spare_reg_activation_13_12;
wire signed[15:0]    spare_reg_activation_13_13;
wire signed[15:0]    spare_reg_activation_13_14;
wire signed[15:0]    spare_reg_activation_13_15;
wire signed[15:0]    spare_reg_activation_13_16;
wire signed[15:0]    spare_reg_activation_13_17;
wire signed[15:0]    spare_reg_activation_13_18;
wire signed[15:0]    spare_reg_activation_13_19;
wire signed[15:0]    spare_reg_activation_13_20;
wire signed[15:0]    spare_reg_activation_13_21;
wire signed[15:0]    spare_reg_activation_13_22;
wire signed[15:0]    spare_reg_activation_13_23;
wire signed[15:0]    spare_reg_activation_13_24;
wire signed[15:0]    spare_reg_activation_13_25;
wire signed[15:0]    spare_reg_activation_13_26;
wire signed[15:0]    spare_reg_activation_13_27;
wire signed[15:0]    spare_reg_activation_13_28;
wire signed[15:0]    spare_reg_activation_13_29;
wire signed[15:0]    spare_reg_activation_13_30;
wire signed[15:0]    spare_reg_activation_13_31;
wire signed[15:0]    spare_reg_activation_14_0;
wire signed[15:0]    spare_reg_activation_14_1;
wire signed[15:0]    spare_reg_activation_14_2;
wire signed[15:0]    spare_reg_activation_14_3;
wire signed[15:0]    spare_reg_activation_14_4;
wire signed[15:0]    spare_reg_activation_14_5;
wire signed[15:0]    spare_reg_activation_14_6;
wire signed[15:0]    spare_reg_activation_14_7;
wire signed[15:0]    spare_reg_activation_14_8;
wire signed[15:0]    spare_reg_activation_14_9;
wire signed[15:0]    spare_reg_activation_14_10;
wire signed[15:0]    spare_reg_activation_14_11;
wire signed[15:0]    spare_reg_activation_14_12;
wire signed[15:0]    spare_reg_activation_14_13;
wire signed[15:0]    spare_reg_activation_14_14;
wire signed[15:0]    spare_reg_activation_14_15;
wire signed[15:0]    spare_reg_activation_14_16;
wire signed[15:0]    spare_reg_activation_14_17;
wire signed[15:0]    spare_reg_activation_14_18;
wire signed[15:0]    spare_reg_activation_14_19;
wire signed[15:0]    spare_reg_activation_14_20;
wire signed[15:0]    spare_reg_activation_14_21;
wire signed[15:0]    spare_reg_activation_14_22;
wire signed[15:0]    spare_reg_activation_14_23;
wire signed[15:0]    spare_reg_activation_14_24;
wire signed[15:0]    spare_reg_activation_14_25;
wire signed[15:0]    spare_reg_activation_14_26;
wire signed[15:0]    spare_reg_activation_14_27;
wire signed[15:0]    spare_reg_activation_14_28;
wire signed[15:0]    spare_reg_activation_14_29;
wire signed[15:0]    spare_reg_activation_14_30;
wire signed[15:0]    spare_reg_activation_14_31;
wire signed[15:0]    spare_reg_activation_15_0;
wire signed[15:0]    spare_reg_activation_15_1;
wire signed[15:0]    spare_reg_activation_15_2;
wire signed[15:0]    spare_reg_activation_15_3;
wire signed[15:0]    spare_reg_activation_15_4;
wire signed[15:0]    spare_reg_activation_15_5;
wire signed[15:0]    spare_reg_activation_15_6;
wire signed[15:0]    spare_reg_activation_15_7;
wire signed[15:0]    spare_reg_activation_15_8;
wire signed[15:0]    spare_reg_activation_15_9;
wire signed[15:0]    spare_reg_activation_15_10;
wire signed[15:0]    spare_reg_activation_15_11;
wire signed[15:0]    spare_reg_activation_15_12;
wire signed[15:0]    spare_reg_activation_15_13;
wire signed[15:0]    spare_reg_activation_15_14;
wire signed[15:0]    spare_reg_activation_15_15;
wire signed[15:0]    spare_reg_activation_15_16;
wire signed[15:0]    spare_reg_activation_15_17;
wire signed[15:0]    spare_reg_activation_15_18;
wire signed[15:0]    spare_reg_activation_15_19;
wire signed[15:0]    spare_reg_activation_15_20;
wire signed[15:0]    spare_reg_activation_15_21;
wire signed[15:0]    spare_reg_activation_15_22;
wire signed[15:0]    spare_reg_activation_15_23;
wire signed[15:0]    spare_reg_activation_15_24;
wire signed[15:0]    spare_reg_activation_15_25;
wire signed[15:0]    spare_reg_activation_15_26;
wire signed[15:0]    spare_reg_activation_15_27;
wire signed[15:0]    spare_reg_activation_15_28;
wire signed[15:0]    spare_reg_activation_15_29;
wire signed[15:0]    spare_reg_activation_15_30;
wire signed[15:0]    spare_reg_activation_15_31;
wire signed[15:0]    spare_reg_activation_16_0;
wire signed[15:0]    spare_reg_activation_16_1;
wire signed[15:0]    spare_reg_activation_16_2;
wire signed[15:0]    spare_reg_activation_16_3;
wire signed[15:0]    spare_reg_activation_16_4;
wire signed[15:0]    spare_reg_activation_16_5;
wire signed[15:0]    spare_reg_activation_16_6;
wire signed[15:0]    spare_reg_activation_16_7;
wire signed[15:0]    spare_reg_activation_16_8;
wire signed[15:0]    spare_reg_activation_16_9;
wire signed[15:0]    spare_reg_activation_16_10;
wire signed[15:0]    spare_reg_activation_16_11;
wire signed[15:0]    spare_reg_activation_16_12;
wire signed[15:0]    spare_reg_activation_16_13;
wire signed[15:0]    spare_reg_activation_16_14;
wire signed[15:0]    spare_reg_activation_16_15;
wire signed[15:0]    spare_reg_activation_16_16;
wire signed[15:0]    spare_reg_activation_16_17;
wire signed[15:0]    spare_reg_activation_16_18;
wire signed[15:0]    spare_reg_activation_16_19;
wire signed[15:0]    spare_reg_activation_16_20;
wire signed[15:0]    spare_reg_activation_16_21;
wire signed[15:0]    spare_reg_activation_16_22;
wire signed[15:0]    spare_reg_activation_16_23;
wire signed[15:0]    spare_reg_activation_16_24;
wire signed[15:0]    spare_reg_activation_16_25;
wire signed[15:0]    spare_reg_activation_16_26;
wire signed[15:0]    spare_reg_activation_16_27;
wire signed[15:0]    spare_reg_activation_16_28;
wire signed[15:0]    spare_reg_activation_16_29;
wire signed[15:0]    spare_reg_activation_16_30;
wire signed[15:0]    spare_reg_activation_16_31;
wire signed[15:0]    spare_reg_activation_17_0;
wire signed[15:0]    spare_reg_activation_17_1;
wire signed[15:0]    spare_reg_activation_17_2;
wire signed[15:0]    spare_reg_activation_17_3;
wire signed[15:0]    spare_reg_activation_17_4;
wire signed[15:0]    spare_reg_activation_17_5;
wire signed[15:0]    spare_reg_activation_17_6;
wire signed[15:0]    spare_reg_activation_17_7;
wire signed[15:0]    spare_reg_activation_17_8;
wire signed[15:0]    spare_reg_activation_17_9;
wire signed[15:0]    spare_reg_activation_17_10;
wire signed[15:0]    spare_reg_activation_17_11;
wire signed[15:0]    spare_reg_activation_17_12;
wire signed[15:0]    spare_reg_activation_17_13;
wire signed[15:0]    spare_reg_activation_17_14;
wire signed[15:0]    spare_reg_activation_17_15;
wire signed[15:0]    spare_reg_activation_17_16;
wire signed[15:0]    spare_reg_activation_17_17;
wire signed[15:0]    spare_reg_activation_17_18;
wire signed[15:0]    spare_reg_activation_17_19;
wire signed[15:0]    spare_reg_activation_17_20;
wire signed[15:0]    spare_reg_activation_17_21;
wire signed[15:0]    spare_reg_activation_17_22;
wire signed[15:0]    spare_reg_activation_17_23;
wire signed[15:0]    spare_reg_activation_17_24;
wire signed[15:0]    spare_reg_activation_17_25;
wire signed[15:0]    spare_reg_activation_17_26;
wire signed[15:0]    spare_reg_activation_17_27;
wire signed[15:0]    spare_reg_activation_17_28;
wire signed[15:0]    spare_reg_activation_17_29;
wire signed[15:0]    spare_reg_activation_17_30;
wire signed[15:0]    spare_reg_activation_17_31;
wire signed[15:0]    spare_reg_activation_18_0;
wire signed[15:0]    spare_reg_activation_18_1;
wire signed[15:0]    spare_reg_activation_18_2;
wire signed[15:0]    spare_reg_activation_18_3;
wire signed[15:0]    spare_reg_activation_18_4;
wire signed[15:0]    spare_reg_activation_18_5;
wire signed[15:0]    spare_reg_activation_18_6;
wire signed[15:0]    spare_reg_activation_18_7;
wire signed[15:0]    spare_reg_activation_18_8;
wire signed[15:0]    spare_reg_activation_18_9;
wire signed[15:0]    spare_reg_activation_18_10;
wire signed[15:0]    spare_reg_activation_18_11;
wire signed[15:0]    spare_reg_activation_18_12;
wire signed[15:0]    spare_reg_activation_18_13;
wire signed[15:0]    spare_reg_activation_18_14;
wire signed[15:0]    spare_reg_activation_18_15;
wire signed[15:0]    spare_reg_activation_18_16;
wire signed[15:0]    spare_reg_activation_18_17;
wire signed[15:0]    spare_reg_activation_18_18;
wire signed[15:0]    spare_reg_activation_18_19;
wire signed[15:0]    spare_reg_activation_18_20;
wire signed[15:0]    spare_reg_activation_18_21;
wire signed[15:0]    spare_reg_activation_18_22;
wire signed[15:0]    spare_reg_activation_18_23;
wire signed[15:0]    spare_reg_activation_18_24;
wire signed[15:0]    spare_reg_activation_18_25;
wire signed[15:0]    spare_reg_activation_18_26;
wire signed[15:0]    spare_reg_activation_18_27;
wire signed[15:0]    spare_reg_activation_18_28;
wire signed[15:0]    spare_reg_activation_18_29;
wire signed[15:0]    spare_reg_activation_18_30;
wire signed[15:0]    spare_reg_activation_18_31;
wire signed[15:0]    spare_reg_activation_19_0;
wire signed[15:0]    spare_reg_activation_19_1;
wire signed[15:0]    spare_reg_activation_19_2;
wire signed[15:0]    spare_reg_activation_19_3;
wire signed[15:0]    spare_reg_activation_19_4;
wire signed[15:0]    spare_reg_activation_19_5;
wire signed[15:0]    spare_reg_activation_19_6;
wire signed[15:0]    spare_reg_activation_19_7;
wire signed[15:0]    spare_reg_activation_19_8;
wire signed[15:0]    spare_reg_activation_19_9;
wire signed[15:0]    spare_reg_activation_19_10;
wire signed[15:0]    spare_reg_activation_19_11;
wire signed[15:0]    spare_reg_activation_19_12;
wire signed[15:0]    spare_reg_activation_19_13;
wire signed[15:0]    spare_reg_activation_19_14;
wire signed[15:0]    spare_reg_activation_19_15;
wire signed[15:0]    spare_reg_activation_19_16;
wire signed[15:0]    spare_reg_activation_19_17;
wire signed[15:0]    spare_reg_activation_19_18;
wire signed[15:0]    spare_reg_activation_19_19;
wire signed[15:0]    spare_reg_activation_19_20;
wire signed[15:0]    spare_reg_activation_19_21;
wire signed[15:0]    spare_reg_activation_19_22;
wire signed[15:0]    spare_reg_activation_19_23;
wire signed[15:0]    spare_reg_activation_19_24;
wire signed[15:0]    spare_reg_activation_19_25;
wire signed[15:0]    spare_reg_activation_19_26;
wire signed[15:0]    spare_reg_activation_19_27;
wire signed[15:0]    spare_reg_activation_19_28;
wire signed[15:0]    spare_reg_activation_19_29;
wire signed[15:0]    spare_reg_activation_19_30;
wire signed[15:0]    spare_reg_activation_19_31;
wire signed[15:0]    spare_reg_activation_20_0;
wire signed[15:0]    spare_reg_activation_20_1;
wire signed[15:0]    spare_reg_activation_20_2;
wire signed[15:0]    spare_reg_activation_20_3;
wire signed[15:0]    spare_reg_activation_20_4;
wire signed[15:0]    spare_reg_activation_20_5;
wire signed[15:0]    spare_reg_activation_20_6;
wire signed[15:0]    spare_reg_activation_20_7;
wire signed[15:0]    spare_reg_activation_20_8;
wire signed[15:0]    spare_reg_activation_20_9;
wire signed[15:0]    spare_reg_activation_20_10;
wire signed[15:0]    spare_reg_activation_20_11;
wire signed[15:0]    spare_reg_activation_20_12;
wire signed[15:0]    spare_reg_activation_20_13;
wire signed[15:0]    spare_reg_activation_20_14;
wire signed[15:0]    spare_reg_activation_20_15;
wire signed[15:0]    spare_reg_activation_20_16;
wire signed[15:0]    spare_reg_activation_20_17;
wire signed[15:0]    spare_reg_activation_20_18;
wire signed[15:0]    spare_reg_activation_20_19;
wire signed[15:0]    spare_reg_activation_20_20;
wire signed[15:0]    spare_reg_activation_20_21;
wire signed[15:0]    spare_reg_activation_20_22;
wire signed[15:0]    spare_reg_activation_20_23;
wire signed[15:0]    spare_reg_activation_20_24;
wire signed[15:0]    spare_reg_activation_20_25;
wire signed[15:0]    spare_reg_activation_20_26;
wire signed[15:0]    spare_reg_activation_20_27;
wire signed[15:0]    spare_reg_activation_20_28;
wire signed[15:0]    spare_reg_activation_20_29;
wire signed[15:0]    spare_reg_activation_20_30;
wire signed[15:0]    spare_reg_activation_20_31;
wire signed[15:0]    spare_reg_activation_21_0;
wire signed[15:0]    spare_reg_activation_21_1;
wire signed[15:0]    spare_reg_activation_21_2;
wire signed[15:0]    spare_reg_activation_21_3;
wire signed[15:0]    spare_reg_activation_21_4;
wire signed[15:0]    spare_reg_activation_21_5;
wire signed[15:0]    spare_reg_activation_21_6;
wire signed[15:0]    spare_reg_activation_21_7;
wire signed[15:0]    spare_reg_activation_21_8;
wire signed[15:0]    spare_reg_activation_21_9;
wire signed[15:0]    spare_reg_activation_21_10;
wire signed[15:0]    spare_reg_activation_21_11;
wire signed[15:0]    spare_reg_activation_21_12;
wire signed[15:0]    spare_reg_activation_21_13;
wire signed[15:0]    spare_reg_activation_21_14;
wire signed[15:0]    spare_reg_activation_21_15;
wire signed[15:0]    spare_reg_activation_21_16;
wire signed[15:0]    spare_reg_activation_21_17;
wire signed[15:0]    spare_reg_activation_21_18;
wire signed[15:0]    spare_reg_activation_21_19;
wire signed[15:0]    spare_reg_activation_21_20;
wire signed[15:0]    spare_reg_activation_21_21;
wire signed[15:0]    spare_reg_activation_21_22;
wire signed[15:0]    spare_reg_activation_21_23;
wire signed[15:0]    spare_reg_activation_21_24;
wire signed[15:0]    spare_reg_activation_21_25;
wire signed[15:0]    spare_reg_activation_21_26;
wire signed[15:0]    spare_reg_activation_21_27;
wire signed[15:0]    spare_reg_activation_21_28;
wire signed[15:0]    spare_reg_activation_21_29;
wire signed[15:0]    spare_reg_activation_21_30;
wire signed[15:0]    spare_reg_activation_21_31;
wire signed[15:0]    spare_reg_activation_22_0;
wire signed[15:0]    spare_reg_activation_22_1;
wire signed[15:0]    spare_reg_activation_22_2;
wire signed[15:0]    spare_reg_activation_22_3;
wire signed[15:0]    spare_reg_activation_22_4;
wire signed[15:0]    spare_reg_activation_22_5;
wire signed[15:0]    spare_reg_activation_22_6;
wire signed[15:0]    spare_reg_activation_22_7;
wire signed[15:0]    spare_reg_activation_22_8;
wire signed[15:0]    spare_reg_activation_22_9;
wire signed[15:0]    spare_reg_activation_22_10;
wire signed[15:0]    spare_reg_activation_22_11;
wire signed[15:0]    spare_reg_activation_22_12;
wire signed[15:0]    spare_reg_activation_22_13;
wire signed[15:0]    spare_reg_activation_22_14;
wire signed[15:0]    spare_reg_activation_22_15;
wire signed[15:0]    spare_reg_activation_22_16;
wire signed[15:0]    spare_reg_activation_22_17;
wire signed[15:0]    spare_reg_activation_22_18;
wire signed[15:0]    spare_reg_activation_22_19;
wire signed[15:0]    spare_reg_activation_22_20;
wire signed[15:0]    spare_reg_activation_22_21;
wire signed[15:0]    spare_reg_activation_22_22;
wire signed[15:0]    spare_reg_activation_22_23;
wire signed[15:0]    spare_reg_activation_22_24;
wire signed[15:0]    spare_reg_activation_22_25;
wire signed[15:0]    spare_reg_activation_22_26;
wire signed[15:0]    spare_reg_activation_22_27;
wire signed[15:0]    spare_reg_activation_22_28;
wire signed[15:0]    spare_reg_activation_22_29;
wire signed[15:0]    spare_reg_activation_22_30;
wire signed[15:0]    spare_reg_activation_22_31;
wire signed[15:0]    spare_reg_activation_23_0;
wire signed[15:0]    spare_reg_activation_23_1;
wire signed[15:0]    spare_reg_activation_23_2;
wire signed[15:0]    spare_reg_activation_23_3;
wire signed[15:0]    spare_reg_activation_23_4;
wire signed[15:0]    spare_reg_activation_23_5;
wire signed[15:0]    spare_reg_activation_23_6;
wire signed[15:0]    spare_reg_activation_23_7;
wire signed[15:0]    spare_reg_activation_23_8;
wire signed[15:0]    spare_reg_activation_23_9;
wire signed[15:0]    spare_reg_activation_23_10;
wire signed[15:0]    spare_reg_activation_23_11;
wire signed[15:0]    spare_reg_activation_23_12;
wire signed[15:0]    spare_reg_activation_23_13;
wire signed[15:0]    spare_reg_activation_23_14;
wire signed[15:0]    spare_reg_activation_23_15;
wire signed[15:0]    spare_reg_activation_23_16;
wire signed[15:0]    spare_reg_activation_23_17;
wire signed[15:0]    spare_reg_activation_23_18;
wire signed[15:0]    spare_reg_activation_23_19;
wire signed[15:0]    spare_reg_activation_23_20;
wire signed[15:0]    spare_reg_activation_23_21;
wire signed[15:0]    spare_reg_activation_23_22;
wire signed[15:0]    spare_reg_activation_23_23;
wire signed[15:0]    spare_reg_activation_23_24;
wire signed[15:0]    spare_reg_activation_23_25;
wire signed[15:0]    spare_reg_activation_23_26;
wire signed[15:0]    spare_reg_activation_23_27;
wire signed[15:0]    spare_reg_activation_23_28;
wire signed[15:0]    spare_reg_activation_23_29;
wire signed[15:0]    spare_reg_activation_23_30;
wire signed[15:0]    spare_reg_activation_23_31;
wire signed[15:0]    spare_reg_activation_24_0;
wire signed[15:0]    spare_reg_activation_24_1;
wire signed[15:0]    spare_reg_activation_24_2;
wire signed[15:0]    spare_reg_activation_24_3;
wire signed[15:0]    spare_reg_activation_24_4;
wire signed[15:0]    spare_reg_activation_24_5;
wire signed[15:0]    spare_reg_activation_24_6;
wire signed[15:0]    spare_reg_activation_24_7;
wire signed[15:0]    spare_reg_activation_24_8;
wire signed[15:0]    spare_reg_activation_24_9;
wire signed[15:0]    spare_reg_activation_24_10;
wire signed[15:0]    spare_reg_activation_24_11;
wire signed[15:0]    spare_reg_activation_24_12;
wire signed[15:0]    spare_reg_activation_24_13;
wire signed[15:0]    spare_reg_activation_24_14;
wire signed[15:0]    spare_reg_activation_24_15;
wire signed[15:0]    spare_reg_activation_24_16;
wire signed[15:0]    spare_reg_activation_24_17;
wire signed[15:0]    spare_reg_activation_24_18;
wire signed[15:0]    spare_reg_activation_24_19;
wire signed[15:0]    spare_reg_activation_24_20;
wire signed[15:0]    spare_reg_activation_24_21;
wire signed[15:0]    spare_reg_activation_24_22;
wire signed[15:0]    spare_reg_activation_24_23;
wire signed[15:0]    spare_reg_activation_24_24;
wire signed[15:0]    spare_reg_activation_24_25;
wire signed[15:0]    spare_reg_activation_24_26;
wire signed[15:0]    spare_reg_activation_24_27;
wire signed[15:0]    spare_reg_activation_24_28;
wire signed[15:0]    spare_reg_activation_24_29;
wire signed[15:0]    spare_reg_activation_24_30;
wire signed[15:0]    spare_reg_activation_24_31;
wire signed[15:0]    spare_reg_activation_25_0;
wire signed[15:0]    spare_reg_activation_25_1;
wire signed[15:0]    spare_reg_activation_25_2;
wire signed[15:0]    spare_reg_activation_25_3;
wire signed[15:0]    spare_reg_activation_25_4;
wire signed[15:0]    spare_reg_activation_25_5;
wire signed[15:0]    spare_reg_activation_25_6;
wire signed[15:0]    spare_reg_activation_25_7;
wire signed[15:0]    spare_reg_activation_25_8;
wire signed[15:0]    spare_reg_activation_25_9;
wire signed[15:0]    spare_reg_activation_25_10;
wire signed[15:0]    spare_reg_activation_25_11;
wire signed[15:0]    spare_reg_activation_25_12;
wire signed[15:0]    spare_reg_activation_25_13;
wire signed[15:0]    spare_reg_activation_25_14;
wire signed[15:0]    spare_reg_activation_25_15;
wire signed[15:0]    spare_reg_activation_25_16;
wire signed[15:0]    spare_reg_activation_25_17;
wire signed[15:0]    spare_reg_activation_25_18;
wire signed[15:0]    spare_reg_activation_25_19;
wire signed[15:0]    spare_reg_activation_25_20;
wire signed[15:0]    spare_reg_activation_25_21;
wire signed[15:0]    spare_reg_activation_25_22;
wire signed[15:0]    spare_reg_activation_25_23;
wire signed[15:0]    spare_reg_activation_25_24;
wire signed[15:0]    spare_reg_activation_25_25;
wire signed[15:0]    spare_reg_activation_25_26;
wire signed[15:0]    spare_reg_activation_25_27;
wire signed[15:0]    spare_reg_activation_25_28;
wire signed[15:0]    spare_reg_activation_25_29;
wire signed[15:0]    spare_reg_activation_25_30;
wire signed[15:0]    spare_reg_activation_25_31;
wire signed[15:0]    spare_reg_activation_26_0;
wire signed[15:0]    spare_reg_activation_26_1;
wire signed[15:0]    spare_reg_activation_26_2;
wire signed[15:0]    spare_reg_activation_26_3;
wire signed[15:0]    spare_reg_activation_26_4;
wire signed[15:0]    spare_reg_activation_26_5;
wire signed[15:0]    spare_reg_activation_26_6;
wire signed[15:0]    spare_reg_activation_26_7;
wire signed[15:0]    spare_reg_activation_26_8;
wire signed[15:0]    spare_reg_activation_26_9;
wire signed[15:0]    spare_reg_activation_26_10;
wire signed[15:0]    spare_reg_activation_26_11;
wire signed[15:0]    spare_reg_activation_26_12;
wire signed[15:0]    spare_reg_activation_26_13;
wire signed[15:0]    spare_reg_activation_26_14;
wire signed[15:0]    spare_reg_activation_26_15;
wire signed[15:0]    spare_reg_activation_26_16;
wire signed[15:0]    spare_reg_activation_26_17;
wire signed[15:0]    spare_reg_activation_26_18;
wire signed[15:0]    spare_reg_activation_26_19;
wire signed[15:0]    spare_reg_activation_26_20;
wire signed[15:0]    spare_reg_activation_26_21;
wire signed[15:0]    spare_reg_activation_26_22;
wire signed[15:0]    spare_reg_activation_26_23;
wire signed[15:0]    spare_reg_activation_26_24;
wire signed[15:0]    spare_reg_activation_26_25;
wire signed[15:0]    spare_reg_activation_26_26;
wire signed[15:0]    spare_reg_activation_26_27;
wire signed[15:0]    spare_reg_activation_26_28;
wire signed[15:0]    spare_reg_activation_26_29;
wire signed[15:0]    spare_reg_activation_26_30;
wire signed[15:0]    spare_reg_activation_26_31;
wire signed[15:0]    spare_reg_activation_27_0;
wire signed[15:0]    spare_reg_activation_27_1;
wire signed[15:0]    spare_reg_activation_27_2;
wire signed[15:0]    spare_reg_activation_27_3;
wire signed[15:0]    spare_reg_activation_27_4;
wire signed[15:0]    spare_reg_activation_27_5;
wire signed[15:0]    spare_reg_activation_27_6;
wire signed[15:0]    spare_reg_activation_27_7;
wire signed[15:0]    spare_reg_activation_27_8;
wire signed[15:0]    spare_reg_activation_27_9;
wire signed[15:0]    spare_reg_activation_27_10;
wire signed[15:0]    spare_reg_activation_27_11;
wire signed[15:0]    spare_reg_activation_27_12;
wire signed[15:0]    spare_reg_activation_27_13;
wire signed[15:0]    spare_reg_activation_27_14;
wire signed[15:0]    spare_reg_activation_27_15;
wire signed[15:0]    spare_reg_activation_27_16;
wire signed[15:0]    spare_reg_activation_27_17;
wire signed[15:0]    spare_reg_activation_27_18;
wire signed[15:0]    spare_reg_activation_27_19;
wire signed[15:0]    spare_reg_activation_27_20;
wire signed[15:0]    spare_reg_activation_27_21;
wire signed[15:0]    spare_reg_activation_27_22;
wire signed[15:0]    spare_reg_activation_27_23;
wire signed[15:0]    spare_reg_activation_27_24;
wire signed[15:0]    spare_reg_activation_27_25;
wire signed[15:0]    spare_reg_activation_27_26;
wire signed[15:0]    spare_reg_activation_27_27;
wire signed[15:0]    spare_reg_activation_27_28;
wire signed[15:0]    spare_reg_activation_27_29;
wire signed[15:0]    spare_reg_activation_27_30;
wire signed[15:0]    spare_reg_activation_27_31;
wire signed[15:0]    spare_reg_activation_28_0;
wire signed[15:0]    spare_reg_activation_28_1;
wire signed[15:0]    spare_reg_activation_28_2;
wire signed[15:0]    spare_reg_activation_28_3;
wire signed[15:0]    spare_reg_activation_28_4;
wire signed[15:0]    spare_reg_activation_28_5;
wire signed[15:0]    spare_reg_activation_28_6;
wire signed[15:0]    spare_reg_activation_28_7;
wire signed[15:0]    spare_reg_activation_28_8;
wire signed[15:0]    spare_reg_activation_28_9;
wire signed[15:0]    spare_reg_activation_28_10;
wire signed[15:0]    spare_reg_activation_28_11;
wire signed[15:0]    spare_reg_activation_28_12;
wire signed[15:0]    spare_reg_activation_28_13;
wire signed[15:0]    spare_reg_activation_28_14;
wire signed[15:0]    spare_reg_activation_28_15;
wire signed[15:0]    spare_reg_activation_28_16;
wire signed[15:0]    spare_reg_activation_28_17;
wire signed[15:0]    spare_reg_activation_28_18;
wire signed[15:0]    spare_reg_activation_28_19;
wire signed[15:0]    spare_reg_activation_28_20;
wire signed[15:0]    spare_reg_activation_28_21;
wire signed[15:0]    spare_reg_activation_28_22;
wire signed[15:0]    spare_reg_activation_28_23;
wire signed[15:0]    spare_reg_activation_28_24;
wire signed[15:0]    spare_reg_activation_28_25;
wire signed[15:0]    spare_reg_activation_28_26;
wire signed[15:0]    spare_reg_activation_28_27;
wire signed[15:0]    spare_reg_activation_28_28;
wire signed[15:0]    spare_reg_activation_28_29;
wire signed[15:0]    spare_reg_activation_28_30;
wire signed[15:0]    spare_reg_activation_28_31;
wire signed[15:0]    spare_reg_activation_29_0;
wire signed[15:0]    spare_reg_activation_29_1;
wire signed[15:0]    spare_reg_activation_29_2;
wire signed[15:0]    spare_reg_activation_29_3;
wire signed[15:0]    spare_reg_activation_29_4;
wire signed[15:0]    spare_reg_activation_29_5;
wire signed[15:0]    spare_reg_activation_29_6;
wire signed[15:0]    spare_reg_activation_29_7;
wire signed[15:0]    spare_reg_activation_29_8;
wire signed[15:0]    spare_reg_activation_29_9;
wire signed[15:0]    spare_reg_activation_29_10;
wire signed[15:0]    spare_reg_activation_29_11;
wire signed[15:0]    spare_reg_activation_29_12;
wire signed[15:0]    spare_reg_activation_29_13;
wire signed[15:0]    spare_reg_activation_29_14;
wire signed[15:0]    spare_reg_activation_29_15;
wire signed[15:0]    spare_reg_activation_29_16;
wire signed[15:0]    spare_reg_activation_29_17;
wire signed[15:0]    spare_reg_activation_29_18;
wire signed[15:0]    spare_reg_activation_29_19;
wire signed[15:0]    spare_reg_activation_29_20;
wire signed[15:0]    spare_reg_activation_29_21;
wire signed[15:0]    spare_reg_activation_29_22;
wire signed[15:0]    spare_reg_activation_29_23;
wire signed[15:0]    spare_reg_activation_29_24;
wire signed[15:0]    spare_reg_activation_29_25;
wire signed[15:0]    spare_reg_activation_29_26;
wire signed[15:0]    spare_reg_activation_29_27;
wire signed[15:0]    spare_reg_activation_29_28;
wire signed[15:0]    spare_reg_activation_29_29;
wire signed[15:0]    spare_reg_activation_29_30;
wire signed[15:0]    spare_reg_activation_29_31;
wire signed[15:0]    spare_reg_activation_30_0;
wire signed[15:0]    spare_reg_activation_30_1;
wire signed[15:0]    spare_reg_activation_30_2;
wire signed[15:0]    spare_reg_activation_30_3;
wire signed[15:0]    spare_reg_activation_30_4;
wire signed[15:0]    spare_reg_activation_30_5;
wire signed[15:0]    spare_reg_activation_30_6;
wire signed[15:0]    spare_reg_activation_30_7;
wire signed[15:0]    spare_reg_activation_30_8;
wire signed[15:0]    spare_reg_activation_30_9;
wire signed[15:0]    spare_reg_activation_30_10;
wire signed[15:0]    spare_reg_activation_30_11;
wire signed[15:0]    spare_reg_activation_30_12;
wire signed[15:0]    spare_reg_activation_30_13;
wire signed[15:0]    spare_reg_activation_30_14;
wire signed[15:0]    spare_reg_activation_30_15;
wire signed[15:0]    spare_reg_activation_30_16;
wire signed[15:0]    spare_reg_activation_30_17;
wire signed[15:0]    spare_reg_activation_30_18;
wire signed[15:0]    spare_reg_activation_30_19;
wire signed[15:0]    spare_reg_activation_30_20;
wire signed[15:0]    spare_reg_activation_30_21;
wire signed[15:0]    spare_reg_activation_30_22;
wire signed[15:0]    spare_reg_activation_30_23;
wire signed[15:0]    spare_reg_activation_30_24;
wire signed[15:0]    spare_reg_activation_30_25;
wire signed[15:0]    spare_reg_activation_30_26;
wire signed[15:0]    spare_reg_activation_30_27;
wire signed[15:0]    spare_reg_activation_30_28;
wire signed[15:0]    spare_reg_activation_30_29;
wire signed[15:0]    spare_reg_activation_30_30;
wire signed[15:0]    spare_reg_activation_30_31;
wire signed[15:0]    spare_reg_activation_31_0;
wire signed[15:0]    spare_reg_activation_31_1;
wire signed[15:0]    spare_reg_activation_31_2;
wire signed[15:0]    spare_reg_activation_31_3;
wire signed[15:0]    spare_reg_activation_31_4;
wire signed[15:0]    spare_reg_activation_31_5;
wire signed[15:0]    spare_reg_activation_31_6;
wire signed[15:0]    spare_reg_activation_31_7;
wire signed[15:0]    spare_reg_activation_31_8;
wire signed[15:0]    spare_reg_activation_31_9;
wire signed[15:0]    spare_reg_activation_31_10;
wire signed[15:0]    spare_reg_activation_31_11;
wire signed[15:0]    spare_reg_activation_31_12;
wire signed[15:0]    spare_reg_activation_31_13;
wire signed[15:0]    spare_reg_activation_31_14;
wire signed[15:0]    spare_reg_activation_31_15;
wire signed[15:0]    spare_reg_activation_31_16;
wire signed[15:0]    spare_reg_activation_31_17;
wire signed[15:0]    spare_reg_activation_31_18;
wire signed[15:0]    spare_reg_activation_31_19;
wire signed[15:0]    spare_reg_activation_31_20;
wire signed[15:0]    spare_reg_activation_31_21;
wire signed[15:0]    spare_reg_activation_31_22;
wire signed[15:0]    spare_reg_activation_31_23;
wire signed[15:0]    spare_reg_activation_31_24;
wire signed[15:0]    spare_reg_activation_31_25;
wire signed[15:0]    spare_reg_activation_31_26;
wire signed[15:0]    spare_reg_activation_31_27;
wire signed[15:0]    spare_reg_activation_31_28;
wire signed[15:0]    spare_reg_activation_31_29;
wire signed[15:0]    spare_reg_activation_31_30;
wire signed[15:0]    spare_reg_activation_31_31;
wire signed[15:0]    spare_reg_weight_0_0;
wire signed[15:0]    spare_reg_psum_0_0;
wire signed[15:0]    spare_reg_weight_0_1;
wire signed[15:0]    spare_reg_psum_0_1;
wire signed[15:0]    spare_reg_weight_0_2;
wire signed[15:0]    spare_reg_psum_0_2;
wire signed[15:0]    spare_reg_weight_0_3;
wire signed[15:0]    spare_reg_psum_0_3;
wire signed[15:0]    spare_reg_weight_0_4;
wire signed[15:0]    spare_reg_psum_0_4;
wire signed[15:0]    spare_reg_weight_0_5;
wire signed[15:0]    spare_reg_psum_0_5;
wire signed[15:0]    spare_reg_weight_0_6;
wire signed[15:0]    spare_reg_psum_0_6;
wire signed[15:0]    spare_reg_weight_0_7;
wire signed[15:0]    spare_reg_psum_0_7;
wire signed[15:0]    spare_reg_weight_0_8;
wire signed[15:0]    spare_reg_psum_0_8;
wire signed[15:0]    spare_reg_weight_0_9;
wire signed[15:0]    spare_reg_psum_0_9;
wire signed[15:0]    spare_reg_weight_0_10;
wire signed[15:0]    spare_reg_psum_0_10;
wire signed[15:0]    spare_reg_weight_0_11;
wire signed[15:0]    spare_reg_psum_0_11;
wire signed[15:0]    spare_reg_weight_0_12;
wire signed[15:0]    spare_reg_psum_0_12;
wire signed[15:0]    spare_reg_weight_0_13;
wire signed[15:0]    spare_reg_psum_0_13;
wire signed[15:0]    spare_reg_weight_0_14;
wire signed[15:0]    spare_reg_psum_0_14;
wire signed[15:0]    spare_reg_weight_0_15;
wire signed[15:0]    spare_reg_psum_0_15;
wire signed[15:0]    spare_reg_weight_0_16;
wire signed[15:0]    spare_reg_psum_0_16;
wire signed[15:0]    spare_reg_weight_0_17;
wire signed[15:0]    spare_reg_psum_0_17;
wire signed[15:0]    spare_reg_weight_0_18;
wire signed[15:0]    spare_reg_psum_0_18;
wire signed[15:0]    spare_reg_weight_0_19;
wire signed[15:0]    spare_reg_psum_0_19;
wire signed[15:0]    spare_reg_weight_0_20;
wire signed[15:0]    spare_reg_psum_0_20;
wire signed[15:0]    spare_reg_weight_0_21;
wire signed[15:0]    spare_reg_psum_0_21;
wire signed[15:0]    spare_reg_weight_0_22;
wire signed[15:0]    spare_reg_psum_0_22;
wire signed[15:0]    spare_reg_weight_0_23;
wire signed[15:0]    spare_reg_psum_0_23;
wire signed[15:0]    spare_reg_weight_0_24;
wire signed[15:0]    spare_reg_psum_0_24;
wire signed[15:0]    spare_reg_weight_0_25;
wire signed[15:0]    spare_reg_psum_0_25;
wire signed[15:0]    spare_reg_weight_0_26;
wire signed[15:0]    spare_reg_psum_0_26;
wire signed[15:0]    spare_reg_weight_0_27;
wire signed[15:0]    spare_reg_psum_0_27;
wire signed[15:0]    spare_reg_weight_0_28;
wire signed[15:0]    spare_reg_psum_0_28;
wire signed[15:0]    spare_reg_weight_0_29;
wire signed[15:0]    spare_reg_psum_0_29;
wire signed[15:0]    spare_reg_weight_0_30;
wire signed[15:0]    spare_reg_psum_0_30;
wire signed[15:0]    spare_reg_weight_0_31;
wire signed[15:0]    spare_reg_psum_0_31;
wire signed[15:0]    spare_reg_weight_1_0;
wire signed[15:0]    spare_reg_psum_1_0;
wire signed[15:0]    spare_reg_weight_1_1;
wire signed[15:0]    spare_reg_psum_1_1;
wire signed[15:0]    spare_reg_weight_1_2;
wire signed[15:0]    spare_reg_psum_1_2;
wire signed[15:0]    spare_reg_weight_1_3;
wire signed[15:0]    spare_reg_psum_1_3;
wire signed[15:0]    spare_reg_weight_1_4;
wire signed[15:0]    spare_reg_psum_1_4;
wire signed[15:0]    spare_reg_weight_1_5;
wire signed[15:0]    spare_reg_psum_1_5;
wire signed[15:0]    spare_reg_weight_1_6;
wire signed[15:0]    spare_reg_psum_1_6;
wire signed[15:0]    spare_reg_weight_1_7;
wire signed[15:0]    spare_reg_psum_1_7;
wire signed[15:0]    spare_reg_weight_1_8;
wire signed[15:0]    spare_reg_psum_1_8;
wire signed[15:0]    spare_reg_weight_1_9;
wire signed[15:0]    spare_reg_psum_1_9;
wire signed[15:0]    spare_reg_weight_1_10;
wire signed[15:0]    spare_reg_psum_1_10;
wire signed[15:0]    spare_reg_weight_1_11;
wire signed[15:0]    spare_reg_psum_1_11;
wire signed[15:0]    spare_reg_weight_1_12;
wire signed[15:0]    spare_reg_psum_1_12;
wire signed[15:0]    spare_reg_weight_1_13;
wire signed[15:0]    spare_reg_psum_1_13;
wire signed[15:0]    spare_reg_weight_1_14;
wire signed[15:0]    spare_reg_psum_1_14;
wire signed[15:0]    spare_reg_weight_1_15;
wire signed[15:0]    spare_reg_psum_1_15;
wire signed[15:0]    spare_reg_weight_1_16;
wire signed[15:0]    spare_reg_psum_1_16;
wire signed[15:0]    spare_reg_weight_1_17;
wire signed[15:0]    spare_reg_psum_1_17;
wire signed[15:0]    spare_reg_weight_1_18;
wire signed[15:0]    spare_reg_psum_1_18;
wire signed[15:0]    spare_reg_weight_1_19;
wire signed[15:0]    spare_reg_psum_1_19;
wire signed[15:0]    spare_reg_weight_1_20;
wire signed[15:0]    spare_reg_psum_1_20;
wire signed[15:0]    spare_reg_weight_1_21;
wire signed[15:0]    spare_reg_psum_1_21;
wire signed[15:0]    spare_reg_weight_1_22;
wire signed[15:0]    spare_reg_psum_1_22;
wire signed[15:0]    spare_reg_weight_1_23;
wire signed[15:0]    spare_reg_psum_1_23;
wire signed[15:0]    spare_reg_weight_1_24;
wire signed[15:0]    spare_reg_psum_1_24;
wire signed[15:0]    spare_reg_weight_1_25;
wire signed[15:0]    spare_reg_psum_1_25;
wire signed[15:0]    spare_reg_weight_1_26;
wire signed[15:0]    spare_reg_psum_1_26;
wire signed[15:0]    spare_reg_weight_1_27;
wire signed[15:0]    spare_reg_psum_1_27;
wire signed[15:0]    spare_reg_weight_1_28;
wire signed[15:0]    spare_reg_psum_1_28;
wire signed[15:0]    spare_reg_weight_1_29;
wire signed[15:0]    spare_reg_psum_1_29;
wire signed[15:0]    spare_reg_weight_1_30;
wire signed[15:0]    spare_reg_psum_1_30;
wire signed[15:0]    spare_reg_weight_1_31;
wire signed[15:0]    spare_reg_psum_1_31;
wire signed[15:0]    spare_reg_weight_2_0;
wire signed[15:0]    spare_reg_psum_2_0;
wire signed[15:0]    spare_reg_weight_2_1;
wire signed[15:0]    spare_reg_psum_2_1;
wire signed[15:0]    spare_reg_weight_2_2;
wire signed[15:0]    spare_reg_psum_2_2;
wire signed[15:0]    spare_reg_weight_2_3;
wire signed[15:0]    spare_reg_psum_2_3;
wire signed[15:0]    spare_reg_weight_2_4;
wire signed[15:0]    spare_reg_psum_2_4;
wire signed[15:0]    spare_reg_weight_2_5;
wire signed[15:0]    spare_reg_psum_2_5;
wire signed[15:0]    spare_reg_weight_2_6;
wire signed[15:0]    spare_reg_psum_2_6;
wire signed[15:0]    spare_reg_weight_2_7;
wire signed[15:0]    spare_reg_psum_2_7;
wire signed[15:0]    spare_reg_weight_2_8;
wire signed[15:0]    spare_reg_psum_2_8;
wire signed[15:0]    spare_reg_weight_2_9;
wire signed[15:0]    spare_reg_psum_2_9;
wire signed[15:0]    spare_reg_weight_2_10;
wire signed[15:0]    spare_reg_psum_2_10;
wire signed[15:0]    spare_reg_weight_2_11;
wire signed[15:0]    spare_reg_psum_2_11;
wire signed[15:0]    spare_reg_weight_2_12;
wire signed[15:0]    spare_reg_psum_2_12;
wire signed[15:0]    spare_reg_weight_2_13;
wire signed[15:0]    spare_reg_psum_2_13;
wire signed[15:0]    spare_reg_weight_2_14;
wire signed[15:0]    spare_reg_psum_2_14;
wire signed[15:0]    spare_reg_weight_2_15;
wire signed[15:0]    spare_reg_psum_2_15;
wire signed[15:0]    spare_reg_weight_2_16;
wire signed[15:0]    spare_reg_psum_2_16;
wire signed[15:0]    spare_reg_weight_2_17;
wire signed[15:0]    spare_reg_psum_2_17;
wire signed[15:0]    spare_reg_weight_2_18;
wire signed[15:0]    spare_reg_psum_2_18;
wire signed[15:0]    spare_reg_weight_2_19;
wire signed[15:0]    spare_reg_psum_2_19;
wire signed[15:0]    spare_reg_weight_2_20;
wire signed[15:0]    spare_reg_psum_2_20;
wire signed[15:0]    spare_reg_weight_2_21;
wire signed[15:0]    spare_reg_psum_2_21;
wire signed[15:0]    spare_reg_weight_2_22;
wire signed[15:0]    spare_reg_psum_2_22;
wire signed[15:0]    spare_reg_weight_2_23;
wire signed[15:0]    spare_reg_psum_2_23;
wire signed[15:0]    spare_reg_weight_2_24;
wire signed[15:0]    spare_reg_psum_2_24;
wire signed[15:0]    spare_reg_weight_2_25;
wire signed[15:0]    spare_reg_psum_2_25;
wire signed[15:0]    spare_reg_weight_2_26;
wire signed[15:0]    spare_reg_psum_2_26;
wire signed[15:0]    spare_reg_weight_2_27;
wire signed[15:0]    spare_reg_psum_2_27;
wire signed[15:0]    spare_reg_weight_2_28;
wire signed[15:0]    spare_reg_psum_2_28;
wire signed[15:0]    spare_reg_weight_2_29;
wire signed[15:0]    spare_reg_psum_2_29;
wire signed[15:0]    spare_reg_weight_2_30;
wire signed[15:0]    spare_reg_psum_2_30;
wire signed[15:0]    spare_reg_weight_2_31;
wire signed[15:0]    spare_reg_psum_2_31;
wire signed[15:0]    spare_reg_weight_3_0;
wire signed[15:0]    spare_reg_psum_3_0;
wire signed[15:0]    spare_reg_weight_3_1;
wire signed[15:0]    spare_reg_psum_3_1;
wire signed[15:0]    spare_reg_weight_3_2;
wire signed[15:0]    spare_reg_psum_3_2;
wire signed[15:0]    spare_reg_weight_3_3;
wire signed[15:0]    spare_reg_psum_3_3;
wire signed[15:0]    spare_reg_weight_3_4;
wire signed[15:0]    spare_reg_psum_3_4;
wire signed[15:0]    spare_reg_weight_3_5;
wire signed[15:0]    spare_reg_psum_3_5;
wire signed[15:0]    spare_reg_weight_3_6;
wire signed[15:0]    spare_reg_psum_3_6;
wire signed[15:0]    spare_reg_weight_3_7;
wire signed[15:0]    spare_reg_psum_3_7;
wire signed[15:0]    spare_reg_weight_3_8;
wire signed[15:0]    spare_reg_psum_3_8;
wire signed[15:0]    spare_reg_weight_3_9;
wire signed[15:0]    spare_reg_psum_3_9;
wire signed[15:0]    spare_reg_weight_3_10;
wire signed[15:0]    spare_reg_psum_3_10;
wire signed[15:0]    spare_reg_weight_3_11;
wire signed[15:0]    spare_reg_psum_3_11;
wire signed[15:0]    spare_reg_weight_3_12;
wire signed[15:0]    spare_reg_psum_3_12;
wire signed[15:0]    spare_reg_weight_3_13;
wire signed[15:0]    spare_reg_psum_3_13;
wire signed[15:0]    spare_reg_weight_3_14;
wire signed[15:0]    spare_reg_psum_3_14;
wire signed[15:0]    spare_reg_weight_3_15;
wire signed[15:0]    spare_reg_psum_3_15;
wire signed[15:0]    spare_reg_weight_3_16;
wire signed[15:0]    spare_reg_psum_3_16;
wire signed[15:0]    spare_reg_weight_3_17;
wire signed[15:0]    spare_reg_psum_3_17;
wire signed[15:0]    spare_reg_weight_3_18;
wire signed[15:0]    spare_reg_psum_3_18;
wire signed[15:0]    spare_reg_weight_3_19;
wire signed[15:0]    spare_reg_psum_3_19;
wire signed[15:0]    spare_reg_weight_3_20;
wire signed[15:0]    spare_reg_psum_3_20;
wire signed[15:0]    spare_reg_weight_3_21;
wire signed[15:0]    spare_reg_psum_3_21;
wire signed[15:0]    spare_reg_weight_3_22;
wire signed[15:0]    spare_reg_psum_3_22;
wire signed[15:0]    spare_reg_weight_3_23;
wire signed[15:0]    spare_reg_psum_3_23;
wire signed[15:0]    spare_reg_weight_3_24;
wire signed[15:0]    spare_reg_psum_3_24;
wire signed[15:0]    spare_reg_weight_3_25;
wire signed[15:0]    spare_reg_psum_3_25;
wire signed[15:0]    spare_reg_weight_3_26;
wire signed[15:0]    spare_reg_psum_3_26;
wire signed[15:0]    spare_reg_weight_3_27;
wire signed[15:0]    spare_reg_psum_3_27;
wire signed[15:0]    spare_reg_weight_3_28;
wire signed[15:0]    spare_reg_psum_3_28;
wire signed[15:0]    spare_reg_weight_3_29;
wire signed[15:0]    spare_reg_psum_3_29;
wire signed[15:0]    spare_reg_weight_3_30;
wire signed[15:0]    spare_reg_psum_3_30;
wire signed[15:0]    spare_reg_weight_3_31;
wire signed[15:0]    spare_reg_psum_3_31;
wire signed[15:0]    spare_reg_weight_4_0;
wire signed[15:0]    spare_reg_psum_4_0;
wire signed[15:0]    spare_reg_weight_4_1;
wire signed[15:0]    spare_reg_psum_4_1;
wire signed[15:0]    spare_reg_weight_4_2;
wire signed[15:0]    spare_reg_psum_4_2;
wire signed[15:0]    spare_reg_weight_4_3;
wire signed[15:0]    spare_reg_psum_4_3;
wire signed[15:0]    spare_reg_weight_4_4;
wire signed[15:0]    spare_reg_psum_4_4;
wire signed[15:0]    spare_reg_weight_4_5;
wire signed[15:0]    spare_reg_psum_4_5;
wire signed[15:0]    spare_reg_weight_4_6;
wire signed[15:0]    spare_reg_psum_4_6;
wire signed[15:0]    spare_reg_weight_4_7;
wire signed[15:0]    spare_reg_psum_4_7;
wire signed[15:0]    spare_reg_weight_4_8;
wire signed[15:0]    spare_reg_psum_4_8;
wire signed[15:0]    spare_reg_weight_4_9;
wire signed[15:0]    spare_reg_psum_4_9;
wire signed[15:0]    spare_reg_weight_4_10;
wire signed[15:0]    spare_reg_psum_4_10;
wire signed[15:0]    spare_reg_weight_4_11;
wire signed[15:0]    spare_reg_psum_4_11;
wire signed[15:0]    spare_reg_weight_4_12;
wire signed[15:0]    spare_reg_psum_4_12;
wire signed[15:0]    spare_reg_weight_4_13;
wire signed[15:0]    spare_reg_psum_4_13;
wire signed[15:0]    spare_reg_weight_4_14;
wire signed[15:0]    spare_reg_psum_4_14;
wire signed[15:0]    spare_reg_weight_4_15;
wire signed[15:0]    spare_reg_psum_4_15;
wire signed[15:0]    spare_reg_weight_4_16;
wire signed[15:0]    spare_reg_psum_4_16;
wire signed[15:0]    spare_reg_weight_4_17;
wire signed[15:0]    spare_reg_psum_4_17;
wire signed[15:0]    spare_reg_weight_4_18;
wire signed[15:0]    spare_reg_psum_4_18;
wire signed[15:0]    spare_reg_weight_4_19;
wire signed[15:0]    spare_reg_psum_4_19;
wire signed[15:0]    spare_reg_weight_4_20;
wire signed[15:0]    spare_reg_psum_4_20;
wire signed[15:0]    spare_reg_weight_4_21;
wire signed[15:0]    spare_reg_psum_4_21;
wire signed[15:0]    spare_reg_weight_4_22;
wire signed[15:0]    spare_reg_psum_4_22;
wire signed[15:0]    spare_reg_weight_4_23;
wire signed[15:0]    spare_reg_psum_4_23;
wire signed[15:0]    spare_reg_weight_4_24;
wire signed[15:0]    spare_reg_psum_4_24;
wire signed[15:0]    spare_reg_weight_4_25;
wire signed[15:0]    spare_reg_psum_4_25;
wire signed[15:0]    spare_reg_weight_4_26;
wire signed[15:0]    spare_reg_psum_4_26;
wire signed[15:0]    spare_reg_weight_4_27;
wire signed[15:0]    spare_reg_psum_4_27;
wire signed[15:0]    spare_reg_weight_4_28;
wire signed[15:0]    spare_reg_psum_4_28;
wire signed[15:0]    spare_reg_weight_4_29;
wire signed[15:0]    spare_reg_psum_4_29;
wire signed[15:0]    spare_reg_weight_4_30;
wire signed[15:0]    spare_reg_psum_4_30;
wire signed[15:0]    spare_reg_weight_4_31;
wire signed[15:0]    spare_reg_psum_4_31;
wire signed[15:0]    spare_reg_weight_5_0;
wire signed[15:0]    spare_reg_psum_5_0;
wire signed[15:0]    spare_reg_weight_5_1;
wire signed[15:0]    spare_reg_psum_5_1;
wire signed[15:0]    spare_reg_weight_5_2;
wire signed[15:0]    spare_reg_psum_5_2;
wire signed[15:0]    spare_reg_weight_5_3;
wire signed[15:0]    spare_reg_psum_5_3;
wire signed[15:0]    spare_reg_weight_5_4;
wire signed[15:0]    spare_reg_psum_5_4;
wire signed[15:0]    spare_reg_weight_5_5;
wire signed[15:0]    spare_reg_psum_5_5;
wire signed[15:0]    spare_reg_weight_5_6;
wire signed[15:0]    spare_reg_psum_5_6;
wire signed[15:0]    spare_reg_weight_5_7;
wire signed[15:0]    spare_reg_psum_5_7;
wire signed[15:0]    spare_reg_weight_5_8;
wire signed[15:0]    spare_reg_psum_5_8;
wire signed[15:0]    spare_reg_weight_5_9;
wire signed[15:0]    spare_reg_psum_5_9;
wire signed[15:0]    spare_reg_weight_5_10;
wire signed[15:0]    spare_reg_psum_5_10;
wire signed[15:0]    spare_reg_weight_5_11;
wire signed[15:0]    spare_reg_psum_5_11;
wire signed[15:0]    spare_reg_weight_5_12;
wire signed[15:0]    spare_reg_psum_5_12;
wire signed[15:0]    spare_reg_weight_5_13;
wire signed[15:0]    spare_reg_psum_5_13;
wire signed[15:0]    spare_reg_weight_5_14;
wire signed[15:0]    spare_reg_psum_5_14;
wire signed[15:0]    spare_reg_weight_5_15;
wire signed[15:0]    spare_reg_psum_5_15;
wire signed[15:0]    spare_reg_weight_5_16;
wire signed[15:0]    spare_reg_psum_5_16;
wire signed[15:0]    spare_reg_weight_5_17;
wire signed[15:0]    spare_reg_psum_5_17;
wire signed[15:0]    spare_reg_weight_5_18;
wire signed[15:0]    spare_reg_psum_5_18;
wire signed[15:0]    spare_reg_weight_5_19;
wire signed[15:0]    spare_reg_psum_5_19;
wire signed[15:0]    spare_reg_weight_5_20;
wire signed[15:0]    spare_reg_psum_5_20;
wire signed[15:0]    spare_reg_weight_5_21;
wire signed[15:0]    spare_reg_psum_5_21;
wire signed[15:0]    spare_reg_weight_5_22;
wire signed[15:0]    spare_reg_psum_5_22;
wire signed[15:0]    spare_reg_weight_5_23;
wire signed[15:0]    spare_reg_psum_5_23;
wire signed[15:0]    spare_reg_weight_5_24;
wire signed[15:0]    spare_reg_psum_5_24;
wire signed[15:0]    spare_reg_weight_5_25;
wire signed[15:0]    spare_reg_psum_5_25;
wire signed[15:0]    spare_reg_weight_5_26;
wire signed[15:0]    spare_reg_psum_5_26;
wire signed[15:0]    spare_reg_weight_5_27;
wire signed[15:0]    spare_reg_psum_5_27;
wire signed[15:0]    spare_reg_weight_5_28;
wire signed[15:0]    spare_reg_psum_5_28;
wire signed[15:0]    spare_reg_weight_5_29;
wire signed[15:0]    spare_reg_psum_5_29;
wire signed[15:0]    spare_reg_weight_5_30;
wire signed[15:0]    spare_reg_psum_5_30;
wire signed[15:0]    spare_reg_weight_5_31;
wire signed[15:0]    spare_reg_psum_5_31;
wire signed[15:0]    spare_reg_weight_6_0;
wire signed[15:0]    spare_reg_psum_6_0;
wire signed[15:0]    spare_reg_weight_6_1;
wire signed[15:0]    spare_reg_psum_6_1;
wire signed[15:0]    spare_reg_weight_6_2;
wire signed[15:0]    spare_reg_psum_6_2;
wire signed[15:0]    spare_reg_weight_6_3;
wire signed[15:0]    spare_reg_psum_6_3;
wire signed[15:0]    spare_reg_weight_6_4;
wire signed[15:0]    spare_reg_psum_6_4;
wire signed[15:0]    spare_reg_weight_6_5;
wire signed[15:0]    spare_reg_psum_6_5;
wire signed[15:0]    spare_reg_weight_6_6;
wire signed[15:0]    spare_reg_psum_6_6;
wire signed[15:0]    spare_reg_weight_6_7;
wire signed[15:0]    spare_reg_psum_6_7;
wire signed[15:0]    spare_reg_weight_6_8;
wire signed[15:0]    spare_reg_psum_6_8;
wire signed[15:0]    spare_reg_weight_6_9;
wire signed[15:0]    spare_reg_psum_6_9;
wire signed[15:0]    spare_reg_weight_6_10;
wire signed[15:0]    spare_reg_psum_6_10;
wire signed[15:0]    spare_reg_weight_6_11;
wire signed[15:0]    spare_reg_psum_6_11;
wire signed[15:0]    spare_reg_weight_6_12;
wire signed[15:0]    spare_reg_psum_6_12;
wire signed[15:0]    spare_reg_weight_6_13;
wire signed[15:0]    spare_reg_psum_6_13;
wire signed[15:0]    spare_reg_weight_6_14;
wire signed[15:0]    spare_reg_psum_6_14;
wire signed[15:0]    spare_reg_weight_6_15;
wire signed[15:0]    spare_reg_psum_6_15;
wire signed[15:0]    spare_reg_weight_6_16;
wire signed[15:0]    spare_reg_psum_6_16;
wire signed[15:0]    spare_reg_weight_6_17;
wire signed[15:0]    spare_reg_psum_6_17;
wire signed[15:0]    spare_reg_weight_6_18;
wire signed[15:0]    spare_reg_psum_6_18;
wire signed[15:0]    spare_reg_weight_6_19;
wire signed[15:0]    spare_reg_psum_6_19;
wire signed[15:0]    spare_reg_weight_6_20;
wire signed[15:0]    spare_reg_psum_6_20;
wire signed[15:0]    spare_reg_weight_6_21;
wire signed[15:0]    spare_reg_psum_6_21;
wire signed[15:0]    spare_reg_weight_6_22;
wire signed[15:0]    spare_reg_psum_6_22;
wire signed[15:0]    spare_reg_weight_6_23;
wire signed[15:0]    spare_reg_psum_6_23;
wire signed[15:0]    spare_reg_weight_6_24;
wire signed[15:0]    spare_reg_psum_6_24;
wire signed[15:0]    spare_reg_weight_6_25;
wire signed[15:0]    spare_reg_psum_6_25;
wire signed[15:0]    spare_reg_weight_6_26;
wire signed[15:0]    spare_reg_psum_6_26;
wire signed[15:0]    spare_reg_weight_6_27;
wire signed[15:0]    spare_reg_psum_6_27;
wire signed[15:0]    spare_reg_weight_6_28;
wire signed[15:0]    spare_reg_psum_6_28;
wire signed[15:0]    spare_reg_weight_6_29;
wire signed[15:0]    spare_reg_psum_6_29;
wire signed[15:0]    spare_reg_weight_6_30;
wire signed[15:0]    spare_reg_psum_6_30;
wire signed[15:0]    spare_reg_weight_6_31;
wire signed[15:0]    spare_reg_psum_6_31;
wire signed[15:0]    spare_reg_weight_7_0;
wire signed[15:0]    spare_reg_psum_7_0;
wire signed[15:0]    spare_reg_weight_7_1;
wire signed[15:0]    spare_reg_psum_7_1;
wire signed[15:0]    spare_reg_weight_7_2;
wire signed[15:0]    spare_reg_psum_7_2;
wire signed[15:0]    spare_reg_weight_7_3;
wire signed[15:0]    spare_reg_psum_7_3;
wire signed[15:0]    spare_reg_weight_7_4;
wire signed[15:0]    spare_reg_psum_7_4;
wire signed[15:0]    spare_reg_weight_7_5;
wire signed[15:0]    spare_reg_psum_7_5;
wire signed[15:0]    spare_reg_weight_7_6;
wire signed[15:0]    spare_reg_psum_7_6;
wire signed[15:0]    spare_reg_weight_7_7;
wire signed[15:0]    spare_reg_psum_7_7;
wire signed[15:0]    spare_reg_weight_7_8;
wire signed[15:0]    spare_reg_psum_7_8;
wire signed[15:0]    spare_reg_weight_7_9;
wire signed[15:0]    spare_reg_psum_7_9;
wire signed[15:0]    spare_reg_weight_7_10;
wire signed[15:0]    spare_reg_psum_7_10;
wire signed[15:0]    spare_reg_weight_7_11;
wire signed[15:0]    spare_reg_psum_7_11;
wire signed[15:0]    spare_reg_weight_7_12;
wire signed[15:0]    spare_reg_psum_7_12;
wire signed[15:0]    spare_reg_weight_7_13;
wire signed[15:0]    spare_reg_psum_7_13;
wire signed[15:0]    spare_reg_weight_7_14;
wire signed[15:0]    spare_reg_psum_7_14;
wire signed[15:0]    spare_reg_weight_7_15;
wire signed[15:0]    spare_reg_psum_7_15;
wire signed[15:0]    spare_reg_weight_7_16;
wire signed[15:0]    spare_reg_psum_7_16;
wire signed[15:0]    spare_reg_weight_7_17;
wire signed[15:0]    spare_reg_psum_7_17;
wire signed[15:0]    spare_reg_weight_7_18;
wire signed[15:0]    spare_reg_psum_7_18;
wire signed[15:0]    spare_reg_weight_7_19;
wire signed[15:0]    spare_reg_psum_7_19;
wire signed[15:0]    spare_reg_weight_7_20;
wire signed[15:0]    spare_reg_psum_7_20;
wire signed[15:0]    spare_reg_weight_7_21;
wire signed[15:0]    spare_reg_psum_7_21;
wire signed[15:0]    spare_reg_weight_7_22;
wire signed[15:0]    spare_reg_psum_7_22;
wire signed[15:0]    spare_reg_weight_7_23;
wire signed[15:0]    spare_reg_psum_7_23;
wire signed[15:0]    spare_reg_weight_7_24;
wire signed[15:0]    spare_reg_psum_7_24;
wire signed[15:0]    spare_reg_weight_7_25;
wire signed[15:0]    spare_reg_psum_7_25;
wire signed[15:0]    spare_reg_weight_7_26;
wire signed[15:0]    spare_reg_psum_7_26;
wire signed[15:0]    spare_reg_weight_7_27;
wire signed[15:0]    spare_reg_psum_7_27;
wire signed[15:0]    spare_reg_weight_7_28;
wire signed[15:0]    spare_reg_psum_7_28;
wire signed[15:0]    spare_reg_weight_7_29;
wire signed[15:0]    spare_reg_psum_7_29;
wire signed[15:0]    spare_reg_weight_7_30;
wire signed[15:0]    spare_reg_psum_7_30;
wire signed[15:0]    spare_reg_weight_7_31;
wire signed[15:0]    spare_reg_psum_7_31;
wire signed[15:0]    spare_reg_weight_8_0;
wire signed[15:0]    spare_reg_psum_8_0;
wire signed[15:0]    spare_reg_weight_8_1;
wire signed[15:0]    spare_reg_psum_8_1;
wire signed[15:0]    spare_reg_weight_8_2;
wire signed[15:0]    spare_reg_psum_8_2;
wire signed[15:0]    spare_reg_weight_8_3;
wire signed[15:0]    spare_reg_psum_8_3;
wire signed[15:0]    spare_reg_weight_8_4;
wire signed[15:0]    spare_reg_psum_8_4;
wire signed[15:0]    spare_reg_weight_8_5;
wire signed[15:0]    spare_reg_psum_8_5;
wire signed[15:0]    spare_reg_weight_8_6;
wire signed[15:0]    spare_reg_psum_8_6;
wire signed[15:0]    spare_reg_weight_8_7;
wire signed[15:0]    spare_reg_psum_8_7;
wire signed[15:0]    spare_reg_weight_8_8;
wire signed[15:0]    spare_reg_psum_8_8;
wire signed[15:0]    spare_reg_weight_8_9;
wire signed[15:0]    spare_reg_psum_8_9;
wire signed[15:0]    spare_reg_weight_8_10;
wire signed[15:0]    spare_reg_psum_8_10;
wire signed[15:0]    spare_reg_weight_8_11;
wire signed[15:0]    spare_reg_psum_8_11;
wire signed[15:0]    spare_reg_weight_8_12;
wire signed[15:0]    spare_reg_psum_8_12;
wire signed[15:0]    spare_reg_weight_8_13;
wire signed[15:0]    spare_reg_psum_8_13;
wire signed[15:0]    spare_reg_weight_8_14;
wire signed[15:0]    spare_reg_psum_8_14;
wire signed[15:0]    spare_reg_weight_8_15;
wire signed[15:0]    spare_reg_psum_8_15;
wire signed[15:0]    spare_reg_weight_8_16;
wire signed[15:0]    spare_reg_psum_8_16;
wire signed[15:0]    spare_reg_weight_8_17;
wire signed[15:0]    spare_reg_psum_8_17;
wire signed[15:0]    spare_reg_weight_8_18;
wire signed[15:0]    spare_reg_psum_8_18;
wire signed[15:0]    spare_reg_weight_8_19;
wire signed[15:0]    spare_reg_psum_8_19;
wire signed[15:0]    spare_reg_weight_8_20;
wire signed[15:0]    spare_reg_psum_8_20;
wire signed[15:0]    spare_reg_weight_8_21;
wire signed[15:0]    spare_reg_psum_8_21;
wire signed[15:0]    spare_reg_weight_8_22;
wire signed[15:0]    spare_reg_psum_8_22;
wire signed[15:0]    spare_reg_weight_8_23;
wire signed[15:0]    spare_reg_psum_8_23;
wire signed[15:0]    spare_reg_weight_8_24;
wire signed[15:0]    spare_reg_psum_8_24;
wire signed[15:0]    spare_reg_weight_8_25;
wire signed[15:0]    spare_reg_psum_8_25;
wire signed[15:0]    spare_reg_weight_8_26;
wire signed[15:0]    spare_reg_psum_8_26;
wire signed[15:0]    spare_reg_weight_8_27;
wire signed[15:0]    spare_reg_psum_8_27;
wire signed[15:0]    spare_reg_weight_8_28;
wire signed[15:0]    spare_reg_psum_8_28;
wire signed[15:0]    spare_reg_weight_8_29;
wire signed[15:0]    spare_reg_psum_8_29;
wire signed[15:0]    spare_reg_weight_8_30;
wire signed[15:0]    spare_reg_psum_8_30;
wire signed[15:0]    spare_reg_weight_8_31;
wire signed[15:0]    spare_reg_psum_8_31;
wire signed[15:0]    spare_reg_weight_9_0;
wire signed[15:0]    spare_reg_psum_9_0;
wire signed[15:0]    spare_reg_weight_9_1;
wire signed[15:0]    spare_reg_psum_9_1;
wire signed[15:0]    spare_reg_weight_9_2;
wire signed[15:0]    spare_reg_psum_9_2;
wire signed[15:0]    spare_reg_weight_9_3;
wire signed[15:0]    spare_reg_psum_9_3;
wire signed[15:0]    spare_reg_weight_9_4;
wire signed[15:0]    spare_reg_psum_9_4;
wire signed[15:0]    spare_reg_weight_9_5;
wire signed[15:0]    spare_reg_psum_9_5;
wire signed[15:0]    spare_reg_weight_9_6;
wire signed[15:0]    spare_reg_psum_9_6;
wire signed[15:0]    spare_reg_weight_9_7;
wire signed[15:0]    spare_reg_psum_9_7;
wire signed[15:0]    spare_reg_weight_9_8;
wire signed[15:0]    spare_reg_psum_9_8;
wire signed[15:0]    spare_reg_weight_9_9;
wire signed[15:0]    spare_reg_psum_9_9;
wire signed[15:0]    spare_reg_weight_9_10;
wire signed[15:0]    spare_reg_psum_9_10;
wire signed[15:0]    spare_reg_weight_9_11;
wire signed[15:0]    spare_reg_psum_9_11;
wire signed[15:0]    spare_reg_weight_9_12;
wire signed[15:0]    spare_reg_psum_9_12;
wire signed[15:0]    spare_reg_weight_9_13;
wire signed[15:0]    spare_reg_psum_9_13;
wire signed[15:0]    spare_reg_weight_9_14;
wire signed[15:0]    spare_reg_psum_9_14;
wire signed[15:0]    spare_reg_weight_9_15;
wire signed[15:0]    spare_reg_psum_9_15;
wire signed[15:0]    spare_reg_weight_9_16;
wire signed[15:0]    spare_reg_psum_9_16;
wire signed[15:0]    spare_reg_weight_9_17;
wire signed[15:0]    spare_reg_psum_9_17;
wire signed[15:0]    spare_reg_weight_9_18;
wire signed[15:0]    spare_reg_psum_9_18;
wire signed[15:0]    spare_reg_weight_9_19;
wire signed[15:0]    spare_reg_psum_9_19;
wire signed[15:0]    spare_reg_weight_9_20;
wire signed[15:0]    spare_reg_psum_9_20;
wire signed[15:0]    spare_reg_weight_9_21;
wire signed[15:0]    spare_reg_psum_9_21;
wire signed[15:0]    spare_reg_weight_9_22;
wire signed[15:0]    spare_reg_psum_9_22;
wire signed[15:0]    spare_reg_weight_9_23;
wire signed[15:0]    spare_reg_psum_9_23;
wire signed[15:0]    spare_reg_weight_9_24;
wire signed[15:0]    spare_reg_psum_9_24;
wire signed[15:0]    spare_reg_weight_9_25;
wire signed[15:0]    spare_reg_psum_9_25;
wire signed[15:0]    spare_reg_weight_9_26;
wire signed[15:0]    spare_reg_psum_9_26;
wire signed[15:0]    spare_reg_weight_9_27;
wire signed[15:0]    spare_reg_psum_9_27;
wire signed[15:0]    spare_reg_weight_9_28;
wire signed[15:0]    spare_reg_psum_9_28;
wire signed[15:0]    spare_reg_weight_9_29;
wire signed[15:0]    spare_reg_psum_9_29;
wire signed[15:0]    spare_reg_weight_9_30;
wire signed[15:0]    spare_reg_psum_9_30;
wire signed[15:0]    spare_reg_weight_9_31;
wire signed[15:0]    spare_reg_psum_9_31;
wire signed[15:0]    spare_reg_weight_10_0;
wire signed[15:0]    spare_reg_psum_10_0;
wire signed[15:0]    spare_reg_weight_10_1;
wire signed[15:0]    spare_reg_psum_10_1;
wire signed[15:0]    spare_reg_weight_10_2;
wire signed[15:0]    spare_reg_psum_10_2;
wire signed[15:0]    spare_reg_weight_10_3;
wire signed[15:0]    spare_reg_psum_10_3;
wire signed[15:0]    spare_reg_weight_10_4;
wire signed[15:0]    spare_reg_psum_10_4;
wire signed[15:0]    spare_reg_weight_10_5;
wire signed[15:0]    spare_reg_psum_10_5;
wire signed[15:0]    spare_reg_weight_10_6;
wire signed[15:0]    spare_reg_psum_10_6;
wire signed[15:0]    spare_reg_weight_10_7;
wire signed[15:0]    spare_reg_psum_10_7;
wire signed[15:0]    spare_reg_weight_10_8;
wire signed[15:0]    spare_reg_psum_10_8;
wire signed[15:0]    spare_reg_weight_10_9;
wire signed[15:0]    spare_reg_psum_10_9;
wire signed[15:0]    spare_reg_weight_10_10;
wire signed[15:0]    spare_reg_psum_10_10;
wire signed[15:0]    spare_reg_weight_10_11;
wire signed[15:0]    spare_reg_psum_10_11;
wire signed[15:0]    spare_reg_weight_10_12;
wire signed[15:0]    spare_reg_psum_10_12;
wire signed[15:0]    spare_reg_weight_10_13;
wire signed[15:0]    spare_reg_psum_10_13;
wire signed[15:0]    spare_reg_weight_10_14;
wire signed[15:0]    spare_reg_psum_10_14;
wire signed[15:0]    spare_reg_weight_10_15;
wire signed[15:0]    spare_reg_psum_10_15;
wire signed[15:0]    spare_reg_weight_10_16;
wire signed[15:0]    spare_reg_psum_10_16;
wire signed[15:0]    spare_reg_weight_10_17;
wire signed[15:0]    spare_reg_psum_10_17;
wire signed[15:0]    spare_reg_weight_10_18;
wire signed[15:0]    spare_reg_psum_10_18;
wire signed[15:0]    spare_reg_weight_10_19;
wire signed[15:0]    spare_reg_psum_10_19;
wire signed[15:0]    spare_reg_weight_10_20;
wire signed[15:0]    spare_reg_psum_10_20;
wire signed[15:0]    spare_reg_weight_10_21;
wire signed[15:0]    spare_reg_psum_10_21;
wire signed[15:0]    spare_reg_weight_10_22;
wire signed[15:0]    spare_reg_psum_10_22;
wire signed[15:0]    spare_reg_weight_10_23;
wire signed[15:0]    spare_reg_psum_10_23;
wire signed[15:0]    spare_reg_weight_10_24;
wire signed[15:0]    spare_reg_psum_10_24;
wire signed[15:0]    spare_reg_weight_10_25;
wire signed[15:0]    spare_reg_psum_10_25;
wire signed[15:0]    spare_reg_weight_10_26;
wire signed[15:0]    spare_reg_psum_10_26;
wire signed[15:0]    spare_reg_weight_10_27;
wire signed[15:0]    spare_reg_psum_10_27;
wire signed[15:0]    spare_reg_weight_10_28;
wire signed[15:0]    spare_reg_psum_10_28;
wire signed[15:0]    spare_reg_weight_10_29;
wire signed[15:0]    spare_reg_psum_10_29;
wire signed[15:0]    spare_reg_weight_10_30;
wire signed[15:0]    spare_reg_psum_10_30;
wire signed[15:0]    spare_reg_weight_10_31;
wire signed[15:0]    spare_reg_psum_10_31;
wire signed[15:0]    spare_reg_weight_11_0;
wire signed[15:0]    spare_reg_psum_11_0;
wire signed[15:0]    spare_reg_weight_11_1;
wire signed[15:0]    spare_reg_psum_11_1;
wire signed[15:0]    spare_reg_weight_11_2;
wire signed[15:0]    spare_reg_psum_11_2;
wire signed[15:0]    spare_reg_weight_11_3;
wire signed[15:0]    spare_reg_psum_11_3;
wire signed[15:0]    spare_reg_weight_11_4;
wire signed[15:0]    spare_reg_psum_11_4;
wire signed[15:0]    spare_reg_weight_11_5;
wire signed[15:0]    spare_reg_psum_11_5;
wire signed[15:0]    spare_reg_weight_11_6;
wire signed[15:0]    spare_reg_psum_11_6;
wire signed[15:0]    spare_reg_weight_11_7;
wire signed[15:0]    spare_reg_psum_11_7;
wire signed[15:0]    spare_reg_weight_11_8;
wire signed[15:0]    spare_reg_psum_11_8;
wire signed[15:0]    spare_reg_weight_11_9;
wire signed[15:0]    spare_reg_psum_11_9;
wire signed[15:0]    spare_reg_weight_11_10;
wire signed[15:0]    spare_reg_psum_11_10;
wire signed[15:0]    spare_reg_weight_11_11;
wire signed[15:0]    spare_reg_psum_11_11;
wire signed[15:0]    spare_reg_weight_11_12;
wire signed[15:0]    spare_reg_psum_11_12;
wire signed[15:0]    spare_reg_weight_11_13;
wire signed[15:0]    spare_reg_psum_11_13;
wire signed[15:0]    spare_reg_weight_11_14;
wire signed[15:0]    spare_reg_psum_11_14;
wire signed[15:0]    spare_reg_weight_11_15;
wire signed[15:0]    spare_reg_psum_11_15;
wire signed[15:0]    spare_reg_weight_11_16;
wire signed[15:0]    spare_reg_psum_11_16;
wire signed[15:0]    spare_reg_weight_11_17;
wire signed[15:0]    spare_reg_psum_11_17;
wire signed[15:0]    spare_reg_weight_11_18;
wire signed[15:0]    spare_reg_psum_11_18;
wire signed[15:0]    spare_reg_weight_11_19;
wire signed[15:0]    spare_reg_psum_11_19;
wire signed[15:0]    spare_reg_weight_11_20;
wire signed[15:0]    spare_reg_psum_11_20;
wire signed[15:0]    spare_reg_weight_11_21;
wire signed[15:0]    spare_reg_psum_11_21;
wire signed[15:0]    spare_reg_weight_11_22;
wire signed[15:0]    spare_reg_psum_11_22;
wire signed[15:0]    spare_reg_weight_11_23;
wire signed[15:0]    spare_reg_psum_11_23;
wire signed[15:0]    spare_reg_weight_11_24;
wire signed[15:0]    spare_reg_psum_11_24;
wire signed[15:0]    spare_reg_weight_11_25;
wire signed[15:0]    spare_reg_psum_11_25;
wire signed[15:0]    spare_reg_weight_11_26;
wire signed[15:0]    spare_reg_psum_11_26;
wire signed[15:0]    spare_reg_weight_11_27;
wire signed[15:0]    spare_reg_psum_11_27;
wire signed[15:0]    spare_reg_weight_11_28;
wire signed[15:0]    spare_reg_psum_11_28;
wire signed[15:0]    spare_reg_weight_11_29;
wire signed[15:0]    spare_reg_psum_11_29;
wire signed[15:0]    spare_reg_weight_11_30;
wire signed[15:0]    spare_reg_psum_11_30;
wire signed[15:0]    spare_reg_weight_11_31;
wire signed[15:0]    spare_reg_psum_11_31;
wire signed[15:0]    spare_reg_weight_12_0;
wire signed[15:0]    spare_reg_psum_12_0;
wire signed[15:0]    spare_reg_weight_12_1;
wire signed[15:0]    spare_reg_psum_12_1;
wire signed[15:0]    spare_reg_weight_12_2;
wire signed[15:0]    spare_reg_psum_12_2;
wire signed[15:0]    spare_reg_weight_12_3;
wire signed[15:0]    spare_reg_psum_12_3;
wire signed[15:0]    spare_reg_weight_12_4;
wire signed[15:0]    spare_reg_psum_12_4;
wire signed[15:0]    spare_reg_weight_12_5;
wire signed[15:0]    spare_reg_psum_12_5;
wire signed[15:0]    spare_reg_weight_12_6;
wire signed[15:0]    spare_reg_psum_12_6;
wire signed[15:0]    spare_reg_weight_12_7;
wire signed[15:0]    spare_reg_psum_12_7;
wire signed[15:0]    spare_reg_weight_12_8;
wire signed[15:0]    spare_reg_psum_12_8;
wire signed[15:0]    spare_reg_weight_12_9;
wire signed[15:0]    spare_reg_psum_12_9;
wire signed[15:0]    spare_reg_weight_12_10;
wire signed[15:0]    spare_reg_psum_12_10;
wire signed[15:0]    spare_reg_weight_12_11;
wire signed[15:0]    spare_reg_psum_12_11;
wire signed[15:0]    spare_reg_weight_12_12;
wire signed[15:0]    spare_reg_psum_12_12;
wire signed[15:0]    spare_reg_weight_12_13;
wire signed[15:0]    spare_reg_psum_12_13;
wire signed[15:0]    spare_reg_weight_12_14;
wire signed[15:0]    spare_reg_psum_12_14;
wire signed[15:0]    spare_reg_weight_12_15;
wire signed[15:0]    spare_reg_psum_12_15;
wire signed[15:0]    spare_reg_weight_12_16;
wire signed[15:0]    spare_reg_psum_12_16;
wire signed[15:0]    spare_reg_weight_12_17;
wire signed[15:0]    spare_reg_psum_12_17;
wire signed[15:0]    spare_reg_weight_12_18;
wire signed[15:0]    spare_reg_psum_12_18;
wire signed[15:0]    spare_reg_weight_12_19;
wire signed[15:0]    spare_reg_psum_12_19;
wire signed[15:0]    spare_reg_weight_12_20;
wire signed[15:0]    spare_reg_psum_12_20;
wire signed[15:0]    spare_reg_weight_12_21;
wire signed[15:0]    spare_reg_psum_12_21;
wire signed[15:0]    spare_reg_weight_12_22;
wire signed[15:0]    spare_reg_psum_12_22;
wire signed[15:0]    spare_reg_weight_12_23;
wire signed[15:0]    spare_reg_psum_12_23;
wire signed[15:0]    spare_reg_weight_12_24;
wire signed[15:0]    spare_reg_psum_12_24;
wire signed[15:0]    spare_reg_weight_12_25;
wire signed[15:0]    spare_reg_psum_12_25;
wire signed[15:0]    spare_reg_weight_12_26;
wire signed[15:0]    spare_reg_psum_12_26;
wire signed[15:0]    spare_reg_weight_12_27;
wire signed[15:0]    spare_reg_psum_12_27;
wire signed[15:0]    spare_reg_weight_12_28;
wire signed[15:0]    spare_reg_psum_12_28;
wire signed[15:0]    spare_reg_weight_12_29;
wire signed[15:0]    spare_reg_psum_12_29;
wire signed[15:0]    spare_reg_weight_12_30;
wire signed[15:0]    spare_reg_psum_12_30;
wire signed[15:0]    spare_reg_weight_12_31;
wire signed[15:0]    spare_reg_psum_12_31;
wire signed[15:0]    spare_reg_weight_13_0;
wire signed[15:0]    spare_reg_psum_13_0;
wire signed[15:0]    spare_reg_weight_13_1;
wire signed[15:0]    spare_reg_psum_13_1;
wire signed[15:0]    spare_reg_weight_13_2;
wire signed[15:0]    spare_reg_psum_13_2;
wire signed[15:0]    spare_reg_weight_13_3;
wire signed[15:0]    spare_reg_psum_13_3;
wire signed[15:0]    spare_reg_weight_13_4;
wire signed[15:0]    spare_reg_psum_13_4;
wire signed[15:0]    spare_reg_weight_13_5;
wire signed[15:0]    spare_reg_psum_13_5;
wire signed[15:0]    spare_reg_weight_13_6;
wire signed[15:0]    spare_reg_psum_13_6;
wire signed[15:0]    spare_reg_weight_13_7;
wire signed[15:0]    spare_reg_psum_13_7;
wire signed[15:0]    spare_reg_weight_13_8;
wire signed[15:0]    spare_reg_psum_13_8;
wire signed[15:0]    spare_reg_weight_13_9;
wire signed[15:0]    spare_reg_psum_13_9;
wire signed[15:0]    spare_reg_weight_13_10;
wire signed[15:0]    spare_reg_psum_13_10;
wire signed[15:0]    spare_reg_weight_13_11;
wire signed[15:0]    spare_reg_psum_13_11;
wire signed[15:0]    spare_reg_weight_13_12;
wire signed[15:0]    spare_reg_psum_13_12;
wire signed[15:0]    spare_reg_weight_13_13;
wire signed[15:0]    spare_reg_psum_13_13;
wire signed[15:0]    spare_reg_weight_13_14;
wire signed[15:0]    spare_reg_psum_13_14;
wire signed[15:0]    spare_reg_weight_13_15;
wire signed[15:0]    spare_reg_psum_13_15;
wire signed[15:0]    spare_reg_weight_13_16;
wire signed[15:0]    spare_reg_psum_13_16;
wire signed[15:0]    spare_reg_weight_13_17;
wire signed[15:0]    spare_reg_psum_13_17;
wire signed[15:0]    spare_reg_weight_13_18;
wire signed[15:0]    spare_reg_psum_13_18;
wire signed[15:0]    spare_reg_weight_13_19;
wire signed[15:0]    spare_reg_psum_13_19;
wire signed[15:0]    spare_reg_weight_13_20;
wire signed[15:0]    spare_reg_psum_13_20;
wire signed[15:0]    spare_reg_weight_13_21;
wire signed[15:0]    spare_reg_psum_13_21;
wire signed[15:0]    spare_reg_weight_13_22;
wire signed[15:0]    spare_reg_psum_13_22;
wire signed[15:0]    spare_reg_weight_13_23;
wire signed[15:0]    spare_reg_psum_13_23;
wire signed[15:0]    spare_reg_weight_13_24;
wire signed[15:0]    spare_reg_psum_13_24;
wire signed[15:0]    spare_reg_weight_13_25;
wire signed[15:0]    spare_reg_psum_13_25;
wire signed[15:0]    spare_reg_weight_13_26;
wire signed[15:0]    spare_reg_psum_13_26;
wire signed[15:0]    spare_reg_weight_13_27;
wire signed[15:0]    spare_reg_psum_13_27;
wire signed[15:0]    spare_reg_weight_13_28;
wire signed[15:0]    spare_reg_psum_13_28;
wire signed[15:0]    spare_reg_weight_13_29;
wire signed[15:0]    spare_reg_psum_13_29;
wire signed[15:0]    spare_reg_weight_13_30;
wire signed[15:0]    spare_reg_psum_13_30;
wire signed[15:0]    spare_reg_weight_13_31;
wire signed[15:0]    spare_reg_psum_13_31;
wire signed[15:0]    spare_reg_weight_14_0;
wire signed[15:0]    spare_reg_psum_14_0;
wire signed[15:0]    spare_reg_weight_14_1;
wire signed[15:0]    spare_reg_psum_14_1;
wire signed[15:0]    spare_reg_weight_14_2;
wire signed[15:0]    spare_reg_psum_14_2;
wire signed[15:0]    spare_reg_weight_14_3;
wire signed[15:0]    spare_reg_psum_14_3;
wire signed[15:0]    spare_reg_weight_14_4;
wire signed[15:0]    spare_reg_psum_14_4;
wire signed[15:0]    spare_reg_weight_14_5;
wire signed[15:0]    spare_reg_psum_14_5;
wire signed[15:0]    spare_reg_weight_14_6;
wire signed[15:0]    spare_reg_psum_14_6;
wire signed[15:0]    spare_reg_weight_14_7;
wire signed[15:0]    spare_reg_psum_14_7;
wire signed[15:0]    spare_reg_weight_14_8;
wire signed[15:0]    spare_reg_psum_14_8;
wire signed[15:0]    spare_reg_weight_14_9;
wire signed[15:0]    spare_reg_psum_14_9;
wire signed[15:0]    spare_reg_weight_14_10;
wire signed[15:0]    spare_reg_psum_14_10;
wire signed[15:0]    spare_reg_weight_14_11;
wire signed[15:0]    spare_reg_psum_14_11;
wire signed[15:0]    spare_reg_weight_14_12;
wire signed[15:0]    spare_reg_psum_14_12;
wire signed[15:0]    spare_reg_weight_14_13;
wire signed[15:0]    spare_reg_psum_14_13;
wire signed[15:0]    spare_reg_weight_14_14;
wire signed[15:0]    spare_reg_psum_14_14;
wire signed[15:0]    spare_reg_weight_14_15;
wire signed[15:0]    spare_reg_psum_14_15;
wire signed[15:0]    spare_reg_weight_14_16;
wire signed[15:0]    spare_reg_psum_14_16;
wire signed[15:0]    spare_reg_weight_14_17;
wire signed[15:0]    spare_reg_psum_14_17;
wire signed[15:0]    spare_reg_weight_14_18;
wire signed[15:0]    spare_reg_psum_14_18;
wire signed[15:0]    spare_reg_weight_14_19;
wire signed[15:0]    spare_reg_psum_14_19;
wire signed[15:0]    spare_reg_weight_14_20;
wire signed[15:0]    spare_reg_psum_14_20;
wire signed[15:0]    spare_reg_weight_14_21;
wire signed[15:0]    spare_reg_psum_14_21;
wire signed[15:0]    spare_reg_weight_14_22;
wire signed[15:0]    spare_reg_psum_14_22;
wire signed[15:0]    spare_reg_weight_14_23;
wire signed[15:0]    spare_reg_psum_14_23;
wire signed[15:0]    spare_reg_weight_14_24;
wire signed[15:0]    spare_reg_psum_14_24;
wire signed[15:0]    spare_reg_weight_14_25;
wire signed[15:0]    spare_reg_psum_14_25;
wire signed[15:0]    spare_reg_weight_14_26;
wire signed[15:0]    spare_reg_psum_14_26;
wire signed[15:0]    spare_reg_weight_14_27;
wire signed[15:0]    spare_reg_psum_14_27;
wire signed[15:0]    spare_reg_weight_14_28;
wire signed[15:0]    spare_reg_psum_14_28;
wire signed[15:0]    spare_reg_weight_14_29;
wire signed[15:0]    spare_reg_psum_14_29;
wire signed[15:0]    spare_reg_weight_14_30;
wire signed[15:0]    spare_reg_psum_14_30;
wire signed[15:0]    spare_reg_weight_14_31;
wire signed[15:0]    spare_reg_psum_14_31;
wire signed[15:0]    spare_reg_weight_15_0;
wire signed[15:0]    spare_reg_psum_15_0;
wire signed[15:0]    spare_reg_weight_15_1;
wire signed[15:0]    spare_reg_psum_15_1;
wire signed[15:0]    spare_reg_weight_15_2;
wire signed[15:0]    spare_reg_psum_15_2;
wire signed[15:0]    spare_reg_weight_15_3;
wire signed[15:0]    spare_reg_psum_15_3;
wire signed[15:0]    spare_reg_weight_15_4;
wire signed[15:0]    spare_reg_psum_15_4;
wire signed[15:0]    spare_reg_weight_15_5;
wire signed[15:0]    spare_reg_psum_15_5;
wire signed[15:0]    spare_reg_weight_15_6;
wire signed[15:0]    spare_reg_psum_15_6;
wire signed[15:0]    spare_reg_weight_15_7;
wire signed[15:0]    spare_reg_psum_15_7;
wire signed[15:0]    spare_reg_weight_15_8;
wire signed[15:0]    spare_reg_psum_15_8;
wire signed[15:0]    spare_reg_weight_15_9;
wire signed[15:0]    spare_reg_psum_15_9;
wire signed[15:0]    spare_reg_weight_15_10;
wire signed[15:0]    spare_reg_psum_15_10;
wire signed[15:0]    spare_reg_weight_15_11;
wire signed[15:0]    spare_reg_psum_15_11;
wire signed[15:0]    spare_reg_weight_15_12;
wire signed[15:0]    spare_reg_psum_15_12;
wire signed[15:0]    spare_reg_weight_15_13;
wire signed[15:0]    spare_reg_psum_15_13;
wire signed[15:0]    spare_reg_weight_15_14;
wire signed[15:0]    spare_reg_psum_15_14;
wire signed[15:0]    spare_reg_weight_15_15;
wire signed[15:0]    spare_reg_psum_15_15;
wire signed[15:0]    spare_reg_weight_15_16;
wire signed[15:0]    spare_reg_psum_15_16;
wire signed[15:0]    spare_reg_weight_15_17;
wire signed[15:0]    spare_reg_psum_15_17;
wire signed[15:0]    spare_reg_weight_15_18;
wire signed[15:0]    spare_reg_psum_15_18;
wire signed[15:0]    spare_reg_weight_15_19;
wire signed[15:0]    spare_reg_psum_15_19;
wire signed[15:0]    spare_reg_weight_15_20;
wire signed[15:0]    spare_reg_psum_15_20;
wire signed[15:0]    spare_reg_weight_15_21;
wire signed[15:0]    spare_reg_psum_15_21;
wire signed[15:0]    spare_reg_weight_15_22;
wire signed[15:0]    spare_reg_psum_15_22;
wire signed[15:0]    spare_reg_weight_15_23;
wire signed[15:0]    spare_reg_psum_15_23;
wire signed[15:0]    spare_reg_weight_15_24;
wire signed[15:0]    spare_reg_psum_15_24;
wire signed[15:0]    spare_reg_weight_15_25;
wire signed[15:0]    spare_reg_psum_15_25;
wire signed[15:0]    spare_reg_weight_15_26;
wire signed[15:0]    spare_reg_psum_15_26;
wire signed[15:0]    spare_reg_weight_15_27;
wire signed[15:0]    spare_reg_psum_15_27;
wire signed[15:0]    spare_reg_weight_15_28;
wire signed[15:0]    spare_reg_psum_15_28;
wire signed[15:0]    spare_reg_weight_15_29;
wire signed[15:0]    spare_reg_psum_15_29;
wire signed[15:0]    spare_reg_weight_15_30;
wire signed[15:0]    spare_reg_psum_15_30;
wire signed[15:0]    spare_reg_weight_15_31;
wire signed[15:0]    spare_reg_psum_15_31;
wire signed[15:0]    spare_reg_weight_16_0;
wire signed[15:0]    spare_reg_psum_16_0;
wire signed[15:0]    spare_reg_weight_16_1;
wire signed[15:0]    spare_reg_psum_16_1;
wire signed[15:0]    spare_reg_weight_16_2;
wire signed[15:0]    spare_reg_psum_16_2;
wire signed[15:0]    spare_reg_weight_16_3;
wire signed[15:0]    spare_reg_psum_16_3;
wire signed[15:0]    spare_reg_weight_16_4;
wire signed[15:0]    spare_reg_psum_16_4;
wire signed[15:0]    spare_reg_weight_16_5;
wire signed[15:0]    spare_reg_psum_16_5;
wire signed[15:0]    spare_reg_weight_16_6;
wire signed[15:0]    spare_reg_psum_16_6;
wire signed[15:0]    spare_reg_weight_16_7;
wire signed[15:0]    spare_reg_psum_16_7;
wire signed[15:0]    spare_reg_weight_16_8;
wire signed[15:0]    spare_reg_psum_16_8;
wire signed[15:0]    spare_reg_weight_16_9;
wire signed[15:0]    spare_reg_psum_16_9;
wire signed[15:0]    spare_reg_weight_16_10;
wire signed[15:0]    spare_reg_psum_16_10;
wire signed[15:0]    spare_reg_weight_16_11;
wire signed[15:0]    spare_reg_psum_16_11;
wire signed[15:0]    spare_reg_weight_16_12;
wire signed[15:0]    spare_reg_psum_16_12;
wire signed[15:0]    spare_reg_weight_16_13;
wire signed[15:0]    spare_reg_psum_16_13;
wire signed[15:0]    spare_reg_weight_16_14;
wire signed[15:0]    spare_reg_psum_16_14;
wire signed[15:0]    spare_reg_weight_16_15;
wire signed[15:0]    spare_reg_psum_16_15;
wire signed[15:0]    spare_reg_weight_16_16;
wire signed[15:0]    spare_reg_psum_16_16;
wire signed[15:0]    spare_reg_weight_16_17;
wire signed[15:0]    spare_reg_psum_16_17;
wire signed[15:0]    spare_reg_weight_16_18;
wire signed[15:0]    spare_reg_psum_16_18;
wire signed[15:0]    spare_reg_weight_16_19;
wire signed[15:0]    spare_reg_psum_16_19;
wire signed[15:0]    spare_reg_weight_16_20;
wire signed[15:0]    spare_reg_psum_16_20;
wire signed[15:0]    spare_reg_weight_16_21;
wire signed[15:0]    spare_reg_psum_16_21;
wire signed[15:0]    spare_reg_weight_16_22;
wire signed[15:0]    spare_reg_psum_16_22;
wire signed[15:0]    spare_reg_weight_16_23;
wire signed[15:0]    spare_reg_psum_16_23;
wire signed[15:0]    spare_reg_weight_16_24;
wire signed[15:0]    spare_reg_psum_16_24;
wire signed[15:0]    spare_reg_weight_16_25;
wire signed[15:0]    spare_reg_psum_16_25;
wire signed[15:0]    spare_reg_weight_16_26;
wire signed[15:0]    spare_reg_psum_16_26;
wire signed[15:0]    spare_reg_weight_16_27;
wire signed[15:0]    spare_reg_psum_16_27;
wire signed[15:0]    spare_reg_weight_16_28;
wire signed[15:0]    spare_reg_psum_16_28;
wire signed[15:0]    spare_reg_weight_16_29;
wire signed[15:0]    spare_reg_psum_16_29;
wire signed[15:0]    spare_reg_weight_16_30;
wire signed[15:0]    spare_reg_psum_16_30;
wire signed[15:0]    spare_reg_weight_16_31;
wire signed[15:0]    spare_reg_psum_16_31;
wire signed[15:0]    spare_reg_weight_17_0;
wire signed[15:0]    spare_reg_psum_17_0;
wire signed[15:0]    spare_reg_weight_17_1;
wire signed[15:0]    spare_reg_psum_17_1;
wire signed[15:0]    spare_reg_weight_17_2;
wire signed[15:0]    spare_reg_psum_17_2;
wire signed[15:0]    spare_reg_weight_17_3;
wire signed[15:0]    spare_reg_psum_17_3;
wire signed[15:0]    spare_reg_weight_17_4;
wire signed[15:0]    spare_reg_psum_17_4;
wire signed[15:0]    spare_reg_weight_17_5;
wire signed[15:0]    spare_reg_psum_17_5;
wire signed[15:0]    spare_reg_weight_17_6;
wire signed[15:0]    spare_reg_psum_17_6;
wire signed[15:0]    spare_reg_weight_17_7;
wire signed[15:0]    spare_reg_psum_17_7;
wire signed[15:0]    spare_reg_weight_17_8;
wire signed[15:0]    spare_reg_psum_17_8;
wire signed[15:0]    spare_reg_weight_17_9;
wire signed[15:0]    spare_reg_psum_17_9;
wire signed[15:0]    spare_reg_weight_17_10;
wire signed[15:0]    spare_reg_psum_17_10;
wire signed[15:0]    spare_reg_weight_17_11;
wire signed[15:0]    spare_reg_psum_17_11;
wire signed[15:0]    spare_reg_weight_17_12;
wire signed[15:0]    spare_reg_psum_17_12;
wire signed[15:0]    spare_reg_weight_17_13;
wire signed[15:0]    spare_reg_psum_17_13;
wire signed[15:0]    spare_reg_weight_17_14;
wire signed[15:0]    spare_reg_psum_17_14;
wire signed[15:0]    spare_reg_weight_17_15;
wire signed[15:0]    spare_reg_psum_17_15;
wire signed[15:0]    spare_reg_weight_17_16;
wire signed[15:0]    spare_reg_psum_17_16;
wire signed[15:0]    spare_reg_weight_17_17;
wire signed[15:0]    spare_reg_psum_17_17;
wire signed[15:0]    spare_reg_weight_17_18;
wire signed[15:0]    spare_reg_psum_17_18;
wire signed[15:0]    spare_reg_weight_17_19;
wire signed[15:0]    spare_reg_psum_17_19;
wire signed[15:0]    spare_reg_weight_17_20;
wire signed[15:0]    spare_reg_psum_17_20;
wire signed[15:0]    spare_reg_weight_17_21;
wire signed[15:0]    spare_reg_psum_17_21;
wire signed[15:0]    spare_reg_weight_17_22;
wire signed[15:0]    spare_reg_psum_17_22;
wire signed[15:0]    spare_reg_weight_17_23;
wire signed[15:0]    spare_reg_psum_17_23;
wire signed[15:0]    spare_reg_weight_17_24;
wire signed[15:0]    spare_reg_psum_17_24;
wire signed[15:0]    spare_reg_weight_17_25;
wire signed[15:0]    spare_reg_psum_17_25;
wire signed[15:0]    spare_reg_weight_17_26;
wire signed[15:0]    spare_reg_psum_17_26;
wire signed[15:0]    spare_reg_weight_17_27;
wire signed[15:0]    spare_reg_psum_17_27;
wire signed[15:0]    spare_reg_weight_17_28;
wire signed[15:0]    spare_reg_psum_17_28;
wire signed[15:0]    spare_reg_weight_17_29;
wire signed[15:0]    spare_reg_psum_17_29;
wire signed[15:0]    spare_reg_weight_17_30;
wire signed[15:0]    spare_reg_psum_17_30;
wire signed[15:0]    spare_reg_weight_17_31;
wire signed[15:0]    spare_reg_psum_17_31;
wire signed[15:0]    spare_reg_weight_18_0;
wire signed[15:0]    spare_reg_psum_18_0;
wire signed[15:0]    spare_reg_weight_18_1;
wire signed[15:0]    spare_reg_psum_18_1;
wire signed[15:0]    spare_reg_weight_18_2;
wire signed[15:0]    spare_reg_psum_18_2;
wire signed[15:0]    spare_reg_weight_18_3;
wire signed[15:0]    spare_reg_psum_18_3;
wire signed[15:0]    spare_reg_weight_18_4;
wire signed[15:0]    spare_reg_psum_18_4;
wire signed[15:0]    spare_reg_weight_18_5;
wire signed[15:0]    spare_reg_psum_18_5;
wire signed[15:0]    spare_reg_weight_18_6;
wire signed[15:0]    spare_reg_psum_18_6;
wire signed[15:0]    spare_reg_weight_18_7;
wire signed[15:0]    spare_reg_psum_18_7;
wire signed[15:0]    spare_reg_weight_18_8;
wire signed[15:0]    spare_reg_psum_18_8;
wire signed[15:0]    spare_reg_weight_18_9;
wire signed[15:0]    spare_reg_psum_18_9;
wire signed[15:0]    spare_reg_weight_18_10;
wire signed[15:0]    spare_reg_psum_18_10;
wire signed[15:0]    spare_reg_weight_18_11;
wire signed[15:0]    spare_reg_psum_18_11;
wire signed[15:0]    spare_reg_weight_18_12;
wire signed[15:0]    spare_reg_psum_18_12;
wire signed[15:0]    spare_reg_weight_18_13;
wire signed[15:0]    spare_reg_psum_18_13;
wire signed[15:0]    spare_reg_weight_18_14;
wire signed[15:0]    spare_reg_psum_18_14;
wire signed[15:0]    spare_reg_weight_18_15;
wire signed[15:0]    spare_reg_psum_18_15;
wire signed[15:0]    spare_reg_weight_18_16;
wire signed[15:0]    spare_reg_psum_18_16;
wire signed[15:0]    spare_reg_weight_18_17;
wire signed[15:0]    spare_reg_psum_18_17;
wire signed[15:0]    spare_reg_weight_18_18;
wire signed[15:0]    spare_reg_psum_18_18;
wire signed[15:0]    spare_reg_weight_18_19;
wire signed[15:0]    spare_reg_psum_18_19;
wire signed[15:0]    spare_reg_weight_18_20;
wire signed[15:0]    spare_reg_psum_18_20;
wire signed[15:0]    spare_reg_weight_18_21;
wire signed[15:0]    spare_reg_psum_18_21;
wire signed[15:0]    spare_reg_weight_18_22;
wire signed[15:0]    spare_reg_psum_18_22;
wire signed[15:0]    spare_reg_weight_18_23;
wire signed[15:0]    spare_reg_psum_18_23;
wire signed[15:0]    spare_reg_weight_18_24;
wire signed[15:0]    spare_reg_psum_18_24;
wire signed[15:0]    spare_reg_weight_18_25;
wire signed[15:0]    spare_reg_psum_18_25;
wire signed[15:0]    spare_reg_weight_18_26;
wire signed[15:0]    spare_reg_psum_18_26;
wire signed[15:0]    spare_reg_weight_18_27;
wire signed[15:0]    spare_reg_psum_18_27;
wire signed[15:0]    spare_reg_weight_18_28;
wire signed[15:0]    spare_reg_psum_18_28;
wire signed[15:0]    spare_reg_weight_18_29;
wire signed[15:0]    spare_reg_psum_18_29;
wire signed[15:0]    spare_reg_weight_18_30;
wire signed[15:0]    spare_reg_psum_18_30;
wire signed[15:0]    spare_reg_weight_18_31;
wire signed[15:0]    spare_reg_psum_18_31;
wire signed[15:0]    spare_reg_weight_19_0;
wire signed[15:0]    spare_reg_psum_19_0;
wire signed[15:0]    spare_reg_weight_19_1;
wire signed[15:0]    spare_reg_psum_19_1;
wire signed[15:0]    spare_reg_weight_19_2;
wire signed[15:0]    spare_reg_psum_19_2;
wire signed[15:0]    spare_reg_weight_19_3;
wire signed[15:0]    spare_reg_psum_19_3;
wire signed[15:0]    spare_reg_weight_19_4;
wire signed[15:0]    spare_reg_psum_19_4;
wire signed[15:0]    spare_reg_weight_19_5;
wire signed[15:0]    spare_reg_psum_19_5;
wire signed[15:0]    spare_reg_weight_19_6;
wire signed[15:0]    spare_reg_psum_19_6;
wire signed[15:0]    spare_reg_weight_19_7;
wire signed[15:0]    spare_reg_psum_19_7;
wire signed[15:0]    spare_reg_weight_19_8;
wire signed[15:0]    spare_reg_psum_19_8;
wire signed[15:0]    spare_reg_weight_19_9;
wire signed[15:0]    spare_reg_psum_19_9;
wire signed[15:0]    spare_reg_weight_19_10;
wire signed[15:0]    spare_reg_psum_19_10;
wire signed[15:0]    spare_reg_weight_19_11;
wire signed[15:0]    spare_reg_psum_19_11;
wire signed[15:0]    spare_reg_weight_19_12;
wire signed[15:0]    spare_reg_psum_19_12;
wire signed[15:0]    spare_reg_weight_19_13;
wire signed[15:0]    spare_reg_psum_19_13;
wire signed[15:0]    spare_reg_weight_19_14;
wire signed[15:0]    spare_reg_psum_19_14;
wire signed[15:0]    spare_reg_weight_19_15;
wire signed[15:0]    spare_reg_psum_19_15;
wire signed[15:0]    spare_reg_weight_19_16;
wire signed[15:0]    spare_reg_psum_19_16;
wire signed[15:0]    spare_reg_weight_19_17;
wire signed[15:0]    spare_reg_psum_19_17;
wire signed[15:0]    spare_reg_weight_19_18;
wire signed[15:0]    spare_reg_psum_19_18;
wire signed[15:0]    spare_reg_weight_19_19;
wire signed[15:0]    spare_reg_psum_19_19;
wire signed[15:0]    spare_reg_weight_19_20;
wire signed[15:0]    spare_reg_psum_19_20;
wire signed[15:0]    spare_reg_weight_19_21;
wire signed[15:0]    spare_reg_psum_19_21;
wire signed[15:0]    spare_reg_weight_19_22;
wire signed[15:0]    spare_reg_psum_19_22;
wire signed[15:0]    spare_reg_weight_19_23;
wire signed[15:0]    spare_reg_psum_19_23;
wire signed[15:0]    spare_reg_weight_19_24;
wire signed[15:0]    spare_reg_psum_19_24;
wire signed[15:0]    spare_reg_weight_19_25;
wire signed[15:0]    spare_reg_psum_19_25;
wire signed[15:0]    spare_reg_weight_19_26;
wire signed[15:0]    spare_reg_psum_19_26;
wire signed[15:0]    spare_reg_weight_19_27;
wire signed[15:0]    spare_reg_psum_19_27;
wire signed[15:0]    spare_reg_weight_19_28;
wire signed[15:0]    spare_reg_psum_19_28;
wire signed[15:0]    spare_reg_weight_19_29;
wire signed[15:0]    spare_reg_psum_19_29;
wire signed[15:0]    spare_reg_weight_19_30;
wire signed[15:0]    spare_reg_psum_19_30;
wire signed[15:0]    spare_reg_weight_19_31;
wire signed[15:0]    spare_reg_psum_19_31;
wire signed[15:0]    spare_reg_weight_20_0;
wire signed[15:0]    spare_reg_psum_20_0;
wire signed[15:0]    spare_reg_weight_20_1;
wire signed[15:0]    spare_reg_psum_20_1;
wire signed[15:0]    spare_reg_weight_20_2;
wire signed[15:0]    spare_reg_psum_20_2;
wire signed[15:0]    spare_reg_weight_20_3;
wire signed[15:0]    spare_reg_psum_20_3;
wire signed[15:0]    spare_reg_weight_20_4;
wire signed[15:0]    spare_reg_psum_20_4;
wire signed[15:0]    spare_reg_weight_20_5;
wire signed[15:0]    spare_reg_psum_20_5;
wire signed[15:0]    spare_reg_weight_20_6;
wire signed[15:0]    spare_reg_psum_20_6;
wire signed[15:0]    spare_reg_weight_20_7;
wire signed[15:0]    spare_reg_psum_20_7;
wire signed[15:0]    spare_reg_weight_20_8;
wire signed[15:0]    spare_reg_psum_20_8;
wire signed[15:0]    spare_reg_weight_20_9;
wire signed[15:0]    spare_reg_psum_20_9;
wire signed[15:0]    spare_reg_weight_20_10;
wire signed[15:0]    spare_reg_psum_20_10;
wire signed[15:0]    spare_reg_weight_20_11;
wire signed[15:0]    spare_reg_psum_20_11;
wire signed[15:0]    spare_reg_weight_20_12;
wire signed[15:0]    spare_reg_psum_20_12;
wire signed[15:0]    spare_reg_weight_20_13;
wire signed[15:0]    spare_reg_psum_20_13;
wire signed[15:0]    spare_reg_weight_20_14;
wire signed[15:0]    spare_reg_psum_20_14;
wire signed[15:0]    spare_reg_weight_20_15;
wire signed[15:0]    spare_reg_psum_20_15;
wire signed[15:0]    spare_reg_weight_20_16;
wire signed[15:0]    spare_reg_psum_20_16;
wire signed[15:0]    spare_reg_weight_20_17;
wire signed[15:0]    spare_reg_psum_20_17;
wire signed[15:0]    spare_reg_weight_20_18;
wire signed[15:0]    spare_reg_psum_20_18;
wire signed[15:0]    spare_reg_weight_20_19;
wire signed[15:0]    spare_reg_psum_20_19;
wire signed[15:0]    spare_reg_weight_20_20;
wire signed[15:0]    spare_reg_psum_20_20;
wire signed[15:0]    spare_reg_weight_20_21;
wire signed[15:0]    spare_reg_psum_20_21;
wire signed[15:0]    spare_reg_weight_20_22;
wire signed[15:0]    spare_reg_psum_20_22;
wire signed[15:0]    spare_reg_weight_20_23;
wire signed[15:0]    spare_reg_psum_20_23;
wire signed[15:0]    spare_reg_weight_20_24;
wire signed[15:0]    spare_reg_psum_20_24;
wire signed[15:0]    spare_reg_weight_20_25;
wire signed[15:0]    spare_reg_psum_20_25;
wire signed[15:0]    spare_reg_weight_20_26;
wire signed[15:0]    spare_reg_psum_20_26;
wire signed[15:0]    spare_reg_weight_20_27;
wire signed[15:0]    spare_reg_psum_20_27;
wire signed[15:0]    spare_reg_weight_20_28;
wire signed[15:0]    spare_reg_psum_20_28;
wire signed[15:0]    spare_reg_weight_20_29;
wire signed[15:0]    spare_reg_psum_20_29;
wire signed[15:0]    spare_reg_weight_20_30;
wire signed[15:0]    spare_reg_psum_20_30;
wire signed[15:0]    spare_reg_weight_20_31;
wire signed[15:0]    spare_reg_psum_20_31;
wire signed[15:0]    spare_reg_weight_21_0;
wire signed[15:0]    spare_reg_psum_21_0;
wire signed[15:0]    spare_reg_weight_21_1;
wire signed[15:0]    spare_reg_psum_21_1;
wire signed[15:0]    spare_reg_weight_21_2;
wire signed[15:0]    spare_reg_psum_21_2;
wire signed[15:0]    spare_reg_weight_21_3;
wire signed[15:0]    spare_reg_psum_21_3;
wire signed[15:0]    spare_reg_weight_21_4;
wire signed[15:0]    spare_reg_psum_21_4;
wire signed[15:0]    spare_reg_weight_21_5;
wire signed[15:0]    spare_reg_psum_21_5;
wire signed[15:0]    spare_reg_weight_21_6;
wire signed[15:0]    spare_reg_psum_21_6;
wire signed[15:0]    spare_reg_weight_21_7;
wire signed[15:0]    spare_reg_psum_21_7;
wire signed[15:0]    spare_reg_weight_21_8;
wire signed[15:0]    spare_reg_psum_21_8;
wire signed[15:0]    spare_reg_weight_21_9;
wire signed[15:0]    spare_reg_psum_21_9;
wire signed[15:0]    spare_reg_weight_21_10;
wire signed[15:0]    spare_reg_psum_21_10;
wire signed[15:0]    spare_reg_weight_21_11;
wire signed[15:0]    spare_reg_psum_21_11;
wire signed[15:0]    spare_reg_weight_21_12;
wire signed[15:0]    spare_reg_psum_21_12;
wire signed[15:0]    spare_reg_weight_21_13;
wire signed[15:0]    spare_reg_psum_21_13;
wire signed[15:0]    spare_reg_weight_21_14;
wire signed[15:0]    spare_reg_psum_21_14;
wire signed[15:0]    spare_reg_weight_21_15;
wire signed[15:0]    spare_reg_psum_21_15;
wire signed[15:0]    spare_reg_weight_21_16;
wire signed[15:0]    spare_reg_psum_21_16;
wire signed[15:0]    spare_reg_weight_21_17;
wire signed[15:0]    spare_reg_psum_21_17;
wire signed[15:0]    spare_reg_weight_21_18;
wire signed[15:0]    spare_reg_psum_21_18;
wire signed[15:0]    spare_reg_weight_21_19;
wire signed[15:0]    spare_reg_psum_21_19;
wire signed[15:0]    spare_reg_weight_21_20;
wire signed[15:0]    spare_reg_psum_21_20;
wire signed[15:0]    spare_reg_weight_21_21;
wire signed[15:0]    spare_reg_psum_21_21;
wire signed[15:0]    spare_reg_weight_21_22;
wire signed[15:0]    spare_reg_psum_21_22;
wire signed[15:0]    spare_reg_weight_21_23;
wire signed[15:0]    spare_reg_psum_21_23;
wire signed[15:0]    spare_reg_weight_21_24;
wire signed[15:0]    spare_reg_psum_21_24;
wire signed[15:0]    spare_reg_weight_21_25;
wire signed[15:0]    spare_reg_psum_21_25;
wire signed[15:0]    spare_reg_weight_21_26;
wire signed[15:0]    spare_reg_psum_21_26;
wire signed[15:0]    spare_reg_weight_21_27;
wire signed[15:0]    spare_reg_psum_21_27;
wire signed[15:0]    spare_reg_weight_21_28;
wire signed[15:0]    spare_reg_psum_21_28;
wire signed[15:0]    spare_reg_weight_21_29;
wire signed[15:0]    spare_reg_psum_21_29;
wire signed[15:0]    spare_reg_weight_21_30;
wire signed[15:0]    spare_reg_psum_21_30;
wire signed[15:0]    spare_reg_weight_21_31;
wire signed[15:0]    spare_reg_psum_21_31;
wire signed[15:0]    spare_reg_weight_22_0;
wire signed[15:0]    spare_reg_psum_22_0;
wire signed[15:0]    spare_reg_weight_22_1;
wire signed[15:0]    spare_reg_psum_22_1;
wire signed[15:0]    spare_reg_weight_22_2;
wire signed[15:0]    spare_reg_psum_22_2;
wire signed[15:0]    spare_reg_weight_22_3;
wire signed[15:0]    spare_reg_psum_22_3;
wire signed[15:0]    spare_reg_weight_22_4;
wire signed[15:0]    spare_reg_psum_22_4;
wire signed[15:0]    spare_reg_weight_22_5;
wire signed[15:0]    spare_reg_psum_22_5;
wire signed[15:0]    spare_reg_weight_22_6;
wire signed[15:0]    spare_reg_psum_22_6;
wire signed[15:0]    spare_reg_weight_22_7;
wire signed[15:0]    spare_reg_psum_22_7;
wire signed[15:0]    spare_reg_weight_22_8;
wire signed[15:0]    spare_reg_psum_22_8;
wire signed[15:0]    spare_reg_weight_22_9;
wire signed[15:0]    spare_reg_psum_22_9;
wire signed[15:0]    spare_reg_weight_22_10;
wire signed[15:0]    spare_reg_psum_22_10;
wire signed[15:0]    spare_reg_weight_22_11;
wire signed[15:0]    spare_reg_psum_22_11;
wire signed[15:0]    spare_reg_weight_22_12;
wire signed[15:0]    spare_reg_psum_22_12;
wire signed[15:0]    spare_reg_weight_22_13;
wire signed[15:0]    spare_reg_psum_22_13;
wire signed[15:0]    spare_reg_weight_22_14;
wire signed[15:0]    spare_reg_psum_22_14;
wire signed[15:0]    spare_reg_weight_22_15;
wire signed[15:0]    spare_reg_psum_22_15;
wire signed[15:0]    spare_reg_weight_22_16;
wire signed[15:0]    spare_reg_psum_22_16;
wire signed[15:0]    spare_reg_weight_22_17;
wire signed[15:0]    spare_reg_psum_22_17;
wire signed[15:0]    spare_reg_weight_22_18;
wire signed[15:0]    spare_reg_psum_22_18;
wire signed[15:0]    spare_reg_weight_22_19;
wire signed[15:0]    spare_reg_psum_22_19;
wire signed[15:0]    spare_reg_weight_22_20;
wire signed[15:0]    spare_reg_psum_22_20;
wire signed[15:0]    spare_reg_weight_22_21;
wire signed[15:0]    spare_reg_psum_22_21;
wire signed[15:0]    spare_reg_weight_22_22;
wire signed[15:0]    spare_reg_psum_22_22;
wire signed[15:0]    spare_reg_weight_22_23;
wire signed[15:0]    spare_reg_psum_22_23;
wire signed[15:0]    spare_reg_weight_22_24;
wire signed[15:0]    spare_reg_psum_22_24;
wire signed[15:0]    spare_reg_weight_22_25;
wire signed[15:0]    spare_reg_psum_22_25;
wire signed[15:0]    spare_reg_weight_22_26;
wire signed[15:0]    spare_reg_psum_22_26;
wire signed[15:0]    spare_reg_weight_22_27;
wire signed[15:0]    spare_reg_psum_22_27;
wire signed[15:0]    spare_reg_weight_22_28;
wire signed[15:0]    spare_reg_psum_22_28;
wire signed[15:0]    spare_reg_weight_22_29;
wire signed[15:0]    spare_reg_psum_22_29;
wire signed[15:0]    spare_reg_weight_22_30;
wire signed[15:0]    spare_reg_psum_22_30;
wire signed[15:0]    spare_reg_weight_22_31;
wire signed[15:0]    spare_reg_psum_22_31;
wire signed[15:0]    spare_reg_weight_23_0;
wire signed[15:0]    spare_reg_psum_23_0;
wire signed[15:0]    spare_reg_weight_23_1;
wire signed[15:0]    spare_reg_psum_23_1;
wire signed[15:0]    spare_reg_weight_23_2;
wire signed[15:0]    spare_reg_psum_23_2;
wire signed[15:0]    spare_reg_weight_23_3;
wire signed[15:0]    spare_reg_psum_23_3;
wire signed[15:0]    spare_reg_weight_23_4;
wire signed[15:0]    spare_reg_psum_23_4;
wire signed[15:0]    spare_reg_weight_23_5;
wire signed[15:0]    spare_reg_psum_23_5;
wire signed[15:0]    spare_reg_weight_23_6;
wire signed[15:0]    spare_reg_psum_23_6;
wire signed[15:0]    spare_reg_weight_23_7;
wire signed[15:0]    spare_reg_psum_23_7;
wire signed[15:0]    spare_reg_weight_23_8;
wire signed[15:0]    spare_reg_psum_23_8;
wire signed[15:0]    spare_reg_weight_23_9;
wire signed[15:0]    spare_reg_psum_23_9;
wire signed[15:0]    spare_reg_weight_23_10;
wire signed[15:0]    spare_reg_psum_23_10;
wire signed[15:0]    spare_reg_weight_23_11;
wire signed[15:0]    spare_reg_psum_23_11;
wire signed[15:0]    spare_reg_weight_23_12;
wire signed[15:0]    spare_reg_psum_23_12;
wire signed[15:0]    spare_reg_weight_23_13;
wire signed[15:0]    spare_reg_psum_23_13;
wire signed[15:0]    spare_reg_weight_23_14;
wire signed[15:0]    spare_reg_psum_23_14;
wire signed[15:0]    spare_reg_weight_23_15;
wire signed[15:0]    spare_reg_psum_23_15;
wire signed[15:0]    spare_reg_weight_23_16;
wire signed[15:0]    spare_reg_psum_23_16;
wire signed[15:0]    spare_reg_weight_23_17;
wire signed[15:0]    spare_reg_psum_23_17;
wire signed[15:0]    spare_reg_weight_23_18;
wire signed[15:0]    spare_reg_psum_23_18;
wire signed[15:0]    spare_reg_weight_23_19;
wire signed[15:0]    spare_reg_psum_23_19;
wire signed[15:0]    spare_reg_weight_23_20;
wire signed[15:0]    spare_reg_psum_23_20;
wire signed[15:0]    spare_reg_weight_23_21;
wire signed[15:0]    spare_reg_psum_23_21;
wire signed[15:0]    spare_reg_weight_23_22;
wire signed[15:0]    spare_reg_psum_23_22;
wire signed[15:0]    spare_reg_weight_23_23;
wire signed[15:0]    spare_reg_psum_23_23;
wire signed[15:0]    spare_reg_weight_23_24;
wire signed[15:0]    spare_reg_psum_23_24;
wire signed[15:0]    spare_reg_weight_23_25;
wire signed[15:0]    spare_reg_psum_23_25;
wire signed[15:0]    spare_reg_weight_23_26;
wire signed[15:0]    spare_reg_psum_23_26;
wire signed[15:0]    spare_reg_weight_23_27;
wire signed[15:0]    spare_reg_psum_23_27;
wire signed[15:0]    spare_reg_weight_23_28;
wire signed[15:0]    spare_reg_psum_23_28;
wire signed[15:0]    spare_reg_weight_23_29;
wire signed[15:0]    spare_reg_psum_23_29;
wire signed[15:0]    spare_reg_weight_23_30;
wire signed[15:0]    spare_reg_psum_23_30;
wire signed[15:0]    spare_reg_weight_23_31;
wire signed[15:0]    spare_reg_psum_23_31;
wire signed[15:0]    spare_reg_weight_24_0;
wire signed[15:0]    spare_reg_psum_24_0;
wire signed[15:0]    spare_reg_weight_24_1;
wire signed[15:0]    spare_reg_psum_24_1;
wire signed[15:0]    spare_reg_weight_24_2;
wire signed[15:0]    spare_reg_psum_24_2;
wire signed[15:0]    spare_reg_weight_24_3;
wire signed[15:0]    spare_reg_psum_24_3;
wire signed[15:0]    spare_reg_weight_24_4;
wire signed[15:0]    spare_reg_psum_24_4;
wire signed[15:0]    spare_reg_weight_24_5;
wire signed[15:0]    spare_reg_psum_24_5;
wire signed[15:0]    spare_reg_weight_24_6;
wire signed[15:0]    spare_reg_psum_24_6;
wire signed[15:0]    spare_reg_weight_24_7;
wire signed[15:0]    spare_reg_psum_24_7;
wire signed[15:0]    spare_reg_weight_24_8;
wire signed[15:0]    spare_reg_psum_24_8;
wire signed[15:0]    spare_reg_weight_24_9;
wire signed[15:0]    spare_reg_psum_24_9;
wire signed[15:0]    spare_reg_weight_24_10;
wire signed[15:0]    spare_reg_psum_24_10;
wire signed[15:0]    spare_reg_weight_24_11;
wire signed[15:0]    spare_reg_psum_24_11;
wire signed[15:0]    spare_reg_weight_24_12;
wire signed[15:0]    spare_reg_psum_24_12;
wire signed[15:0]    spare_reg_weight_24_13;
wire signed[15:0]    spare_reg_psum_24_13;
wire signed[15:0]    spare_reg_weight_24_14;
wire signed[15:0]    spare_reg_psum_24_14;
wire signed[15:0]    spare_reg_weight_24_15;
wire signed[15:0]    spare_reg_psum_24_15;
wire signed[15:0]    spare_reg_weight_24_16;
wire signed[15:0]    spare_reg_psum_24_16;
wire signed[15:0]    spare_reg_weight_24_17;
wire signed[15:0]    spare_reg_psum_24_17;
wire signed[15:0]    spare_reg_weight_24_18;
wire signed[15:0]    spare_reg_psum_24_18;
wire signed[15:0]    spare_reg_weight_24_19;
wire signed[15:0]    spare_reg_psum_24_19;
wire signed[15:0]    spare_reg_weight_24_20;
wire signed[15:0]    spare_reg_psum_24_20;
wire signed[15:0]    spare_reg_weight_24_21;
wire signed[15:0]    spare_reg_psum_24_21;
wire signed[15:0]    spare_reg_weight_24_22;
wire signed[15:0]    spare_reg_psum_24_22;
wire signed[15:0]    spare_reg_weight_24_23;
wire signed[15:0]    spare_reg_psum_24_23;
wire signed[15:0]    spare_reg_weight_24_24;
wire signed[15:0]    spare_reg_psum_24_24;
wire signed[15:0]    spare_reg_weight_24_25;
wire signed[15:0]    spare_reg_psum_24_25;
wire signed[15:0]    spare_reg_weight_24_26;
wire signed[15:0]    spare_reg_psum_24_26;
wire signed[15:0]    spare_reg_weight_24_27;
wire signed[15:0]    spare_reg_psum_24_27;
wire signed[15:0]    spare_reg_weight_24_28;
wire signed[15:0]    spare_reg_psum_24_28;
wire signed[15:0]    spare_reg_weight_24_29;
wire signed[15:0]    spare_reg_psum_24_29;
wire signed[15:0]    spare_reg_weight_24_30;
wire signed[15:0]    spare_reg_psum_24_30;
wire signed[15:0]    spare_reg_weight_24_31;
wire signed[15:0]    spare_reg_psum_24_31;
wire signed[15:0]    spare_reg_weight_25_0;
wire signed[15:0]    spare_reg_psum_25_0;
wire signed[15:0]    spare_reg_weight_25_1;
wire signed[15:0]    spare_reg_psum_25_1;
wire signed[15:0]    spare_reg_weight_25_2;
wire signed[15:0]    spare_reg_psum_25_2;
wire signed[15:0]    spare_reg_weight_25_3;
wire signed[15:0]    spare_reg_psum_25_3;
wire signed[15:0]    spare_reg_weight_25_4;
wire signed[15:0]    spare_reg_psum_25_4;
wire signed[15:0]    spare_reg_weight_25_5;
wire signed[15:0]    spare_reg_psum_25_5;
wire signed[15:0]    spare_reg_weight_25_6;
wire signed[15:0]    spare_reg_psum_25_6;
wire signed[15:0]    spare_reg_weight_25_7;
wire signed[15:0]    spare_reg_psum_25_7;
wire signed[15:0]    spare_reg_weight_25_8;
wire signed[15:0]    spare_reg_psum_25_8;
wire signed[15:0]    spare_reg_weight_25_9;
wire signed[15:0]    spare_reg_psum_25_9;
wire signed[15:0]    spare_reg_weight_25_10;
wire signed[15:0]    spare_reg_psum_25_10;
wire signed[15:0]    spare_reg_weight_25_11;
wire signed[15:0]    spare_reg_psum_25_11;
wire signed[15:0]    spare_reg_weight_25_12;
wire signed[15:0]    spare_reg_psum_25_12;
wire signed[15:0]    spare_reg_weight_25_13;
wire signed[15:0]    spare_reg_psum_25_13;
wire signed[15:0]    spare_reg_weight_25_14;
wire signed[15:0]    spare_reg_psum_25_14;
wire signed[15:0]    spare_reg_weight_25_15;
wire signed[15:0]    spare_reg_psum_25_15;
wire signed[15:0]    spare_reg_weight_25_16;
wire signed[15:0]    spare_reg_psum_25_16;
wire signed[15:0]    spare_reg_weight_25_17;
wire signed[15:0]    spare_reg_psum_25_17;
wire signed[15:0]    spare_reg_weight_25_18;
wire signed[15:0]    spare_reg_psum_25_18;
wire signed[15:0]    spare_reg_weight_25_19;
wire signed[15:0]    spare_reg_psum_25_19;
wire signed[15:0]    spare_reg_weight_25_20;
wire signed[15:0]    spare_reg_psum_25_20;
wire signed[15:0]    spare_reg_weight_25_21;
wire signed[15:0]    spare_reg_psum_25_21;
wire signed[15:0]    spare_reg_weight_25_22;
wire signed[15:0]    spare_reg_psum_25_22;
wire signed[15:0]    spare_reg_weight_25_23;
wire signed[15:0]    spare_reg_psum_25_23;
wire signed[15:0]    spare_reg_weight_25_24;
wire signed[15:0]    spare_reg_psum_25_24;
wire signed[15:0]    spare_reg_weight_25_25;
wire signed[15:0]    spare_reg_psum_25_25;
wire signed[15:0]    spare_reg_weight_25_26;
wire signed[15:0]    spare_reg_psum_25_26;
wire signed[15:0]    spare_reg_weight_25_27;
wire signed[15:0]    spare_reg_psum_25_27;
wire signed[15:0]    spare_reg_weight_25_28;
wire signed[15:0]    spare_reg_psum_25_28;
wire signed[15:0]    spare_reg_weight_25_29;
wire signed[15:0]    spare_reg_psum_25_29;
wire signed[15:0]    spare_reg_weight_25_30;
wire signed[15:0]    spare_reg_psum_25_30;
wire signed[15:0]    spare_reg_weight_25_31;
wire signed[15:0]    spare_reg_psum_25_31;
wire signed[15:0]    spare_reg_weight_26_0;
wire signed[15:0]    spare_reg_psum_26_0;
wire signed[15:0]    spare_reg_weight_26_1;
wire signed[15:0]    spare_reg_psum_26_1;
wire signed[15:0]    spare_reg_weight_26_2;
wire signed[15:0]    spare_reg_psum_26_2;
wire signed[15:0]    spare_reg_weight_26_3;
wire signed[15:0]    spare_reg_psum_26_3;
wire signed[15:0]    spare_reg_weight_26_4;
wire signed[15:0]    spare_reg_psum_26_4;
wire signed[15:0]    spare_reg_weight_26_5;
wire signed[15:0]    spare_reg_psum_26_5;
wire signed[15:0]    spare_reg_weight_26_6;
wire signed[15:0]    spare_reg_psum_26_6;
wire signed[15:0]    spare_reg_weight_26_7;
wire signed[15:0]    spare_reg_psum_26_7;
wire signed[15:0]    spare_reg_weight_26_8;
wire signed[15:0]    spare_reg_psum_26_8;
wire signed[15:0]    spare_reg_weight_26_9;
wire signed[15:0]    spare_reg_psum_26_9;
wire signed[15:0]    spare_reg_weight_26_10;
wire signed[15:0]    spare_reg_psum_26_10;
wire signed[15:0]    spare_reg_weight_26_11;
wire signed[15:0]    spare_reg_psum_26_11;
wire signed[15:0]    spare_reg_weight_26_12;
wire signed[15:0]    spare_reg_psum_26_12;
wire signed[15:0]    spare_reg_weight_26_13;
wire signed[15:0]    spare_reg_psum_26_13;
wire signed[15:0]    spare_reg_weight_26_14;
wire signed[15:0]    spare_reg_psum_26_14;
wire signed[15:0]    spare_reg_weight_26_15;
wire signed[15:0]    spare_reg_psum_26_15;
wire signed[15:0]    spare_reg_weight_26_16;
wire signed[15:0]    spare_reg_psum_26_16;
wire signed[15:0]    spare_reg_weight_26_17;
wire signed[15:0]    spare_reg_psum_26_17;
wire signed[15:0]    spare_reg_weight_26_18;
wire signed[15:0]    spare_reg_psum_26_18;
wire signed[15:0]    spare_reg_weight_26_19;
wire signed[15:0]    spare_reg_psum_26_19;
wire signed[15:0]    spare_reg_weight_26_20;
wire signed[15:0]    spare_reg_psum_26_20;
wire signed[15:0]    spare_reg_weight_26_21;
wire signed[15:0]    spare_reg_psum_26_21;
wire signed[15:0]    spare_reg_weight_26_22;
wire signed[15:0]    spare_reg_psum_26_22;
wire signed[15:0]    spare_reg_weight_26_23;
wire signed[15:0]    spare_reg_psum_26_23;
wire signed[15:0]    spare_reg_weight_26_24;
wire signed[15:0]    spare_reg_psum_26_24;
wire signed[15:0]    spare_reg_weight_26_25;
wire signed[15:0]    spare_reg_psum_26_25;
wire signed[15:0]    spare_reg_weight_26_26;
wire signed[15:0]    spare_reg_psum_26_26;
wire signed[15:0]    spare_reg_weight_26_27;
wire signed[15:0]    spare_reg_psum_26_27;
wire signed[15:0]    spare_reg_weight_26_28;
wire signed[15:0]    spare_reg_psum_26_28;
wire signed[15:0]    spare_reg_weight_26_29;
wire signed[15:0]    spare_reg_psum_26_29;
wire signed[15:0]    spare_reg_weight_26_30;
wire signed[15:0]    spare_reg_psum_26_30;
wire signed[15:0]    spare_reg_weight_26_31;
wire signed[15:0]    spare_reg_psum_26_31;
wire signed[15:0]    spare_reg_weight_27_0;
wire signed[15:0]    spare_reg_psum_27_0;
wire signed[15:0]    spare_reg_weight_27_1;
wire signed[15:0]    spare_reg_psum_27_1;
wire signed[15:0]    spare_reg_weight_27_2;
wire signed[15:0]    spare_reg_psum_27_2;
wire signed[15:0]    spare_reg_weight_27_3;
wire signed[15:0]    spare_reg_psum_27_3;
wire signed[15:0]    spare_reg_weight_27_4;
wire signed[15:0]    spare_reg_psum_27_4;
wire signed[15:0]    spare_reg_weight_27_5;
wire signed[15:0]    spare_reg_psum_27_5;
wire signed[15:0]    spare_reg_weight_27_6;
wire signed[15:0]    spare_reg_psum_27_6;
wire signed[15:0]    spare_reg_weight_27_7;
wire signed[15:0]    spare_reg_psum_27_7;
wire signed[15:0]    spare_reg_weight_27_8;
wire signed[15:0]    spare_reg_psum_27_8;
wire signed[15:0]    spare_reg_weight_27_9;
wire signed[15:0]    spare_reg_psum_27_9;
wire signed[15:0]    spare_reg_weight_27_10;
wire signed[15:0]    spare_reg_psum_27_10;
wire signed[15:0]    spare_reg_weight_27_11;
wire signed[15:0]    spare_reg_psum_27_11;
wire signed[15:0]    spare_reg_weight_27_12;
wire signed[15:0]    spare_reg_psum_27_12;
wire signed[15:0]    spare_reg_weight_27_13;
wire signed[15:0]    spare_reg_psum_27_13;
wire signed[15:0]    spare_reg_weight_27_14;
wire signed[15:0]    spare_reg_psum_27_14;
wire signed[15:0]    spare_reg_weight_27_15;
wire signed[15:0]    spare_reg_psum_27_15;
wire signed[15:0]    spare_reg_weight_27_16;
wire signed[15:0]    spare_reg_psum_27_16;
wire signed[15:0]    spare_reg_weight_27_17;
wire signed[15:0]    spare_reg_psum_27_17;
wire signed[15:0]    spare_reg_weight_27_18;
wire signed[15:0]    spare_reg_psum_27_18;
wire signed[15:0]    spare_reg_weight_27_19;
wire signed[15:0]    spare_reg_psum_27_19;
wire signed[15:0]    spare_reg_weight_27_20;
wire signed[15:0]    spare_reg_psum_27_20;
wire signed[15:0]    spare_reg_weight_27_21;
wire signed[15:0]    spare_reg_psum_27_21;
wire signed[15:0]    spare_reg_weight_27_22;
wire signed[15:0]    spare_reg_psum_27_22;
wire signed[15:0]    spare_reg_weight_27_23;
wire signed[15:0]    spare_reg_psum_27_23;
wire signed[15:0]    spare_reg_weight_27_24;
wire signed[15:0]    spare_reg_psum_27_24;
wire signed[15:0]    spare_reg_weight_27_25;
wire signed[15:0]    spare_reg_psum_27_25;
wire signed[15:0]    spare_reg_weight_27_26;
wire signed[15:0]    spare_reg_psum_27_26;
wire signed[15:0]    spare_reg_weight_27_27;
wire signed[15:0]    spare_reg_psum_27_27;
wire signed[15:0]    spare_reg_weight_27_28;
wire signed[15:0]    spare_reg_psum_27_28;
wire signed[15:0]    spare_reg_weight_27_29;
wire signed[15:0]    spare_reg_psum_27_29;
wire signed[15:0]    spare_reg_weight_27_30;
wire signed[15:0]    spare_reg_psum_27_30;
wire signed[15:0]    spare_reg_weight_27_31;
wire signed[15:0]    spare_reg_psum_27_31;
wire signed[15:0]    spare_reg_weight_28_0;
wire signed[15:0]    spare_reg_psum_28_0;
wire signed[15:0]    spare_reg_weight_28_1;
wire signed[15:0]    spare_reg_psum_28_1;
wire signed[15:0]    spare_reg_weight_28_2;
wire signed[15:0]    spare_reg_psum_28_2;
wire signed[15:0]    spare_reg_weight_28_3;
wire signed[15:0]    spare_reg_psum_28_3;
wire signed[15:0]    spare_reg_weight_28_4;
wire signed[15:0]    spare_reg_psum_28_4;
wire signed[15:0]    spare_reg_weight_28_5;
wire signed[15:0]    spare_reg_psum_28_5;
wire signed[15:0]    spare_reg_weight_28_6;
wire signed[15:0]    spare_reg_psum_28_6;
wire signed[15:0]    spare_reg_weight_28_7;
wire signed[15:0]    spare_reg_psum_28_7;
wire signed[15:0]    spare_reg_weight_28_8;
wire signed[15:0]    spare_reg_psum_28_8;
wire signed[15:0]    spare_reg_weight_28_9;
wire signed[15:0]    spare_reg_psum_28_9;
wire signed[15:0]    spare_reg_weight_28_10;
wire signed[15:0]    spare_reg_psum_28_10;
wire signed[15:0]    spare_reg_weight_28_11;
wire signed[15:0]    spare_reg_psum_28_11;
wire signed[15:0]    spare_reg_weight_28_12;
wire signed[15:0]    spare_reg_psum_28_12;
wire signed[15:0]    spare_reg_weight_28_13;
wire signed[15:0]    spare_reg_psum_28_13;
wire signed[15:0]    spare_reg_weight_28_14;
wire signed[15:0]    spare_reg_psum_28_14;
wire signed[15:0]    spare_reg_weight_28_15;
wire signed[15:0]    spare_reg_psum_28_15;
wire signed[15:0]    spare_reg_weight_28_16;
wire signed[15:0]    spare_reg_psum_28_16;
wire signed[15:0]    spare_reg_weight_28_17;
wire signed[15:0]    spare_reg_psum_28_17;
wire signed[15:0]    spare_reg_weight_28_18;
wire signed[15:0]    spare_reg_psum_28_18;
wire signed[15:0]    spare_reg_weight_28_19;
wire signed[15:0]    spare_reg_psum_28_19;
wire signed[15:0]    spare_reg_weight_28_20;
wire signed[15:0]    spare_reg_psum_28_20;
wire signed[15:0]    spare_reg_weight_28_21;
wire signed[15:0]    spare_reg_psum_28_21;
wire signed[15:0]    spare_reg_weight_28_22;
wire signed[15:0]    spare_reg_psum_28_22;
wire signed[15:0]    spare_reg_weight_28_23;
wire signed[15:0]    spare_reg_psum_28_23;
wire signed[15:0]    spare_reg_weight_28_24;
wire signed[15:0]    spare_reg_psum_28_24;
wire signed[15:0]    spare_reg_weight_28_25;
wire signed[15:0]    spare_reg_psum_28_25;
wire signed[15:0]    spare_reg_weight_28_26;
wire signed[15:0]    spare_reg_psum_28_26;
wire signed[15:0]    spare_reg_weight_28_27;
wire signed[15:0]    spare_reg_psum_28_27;
wire signed[15:0]    spare_reg_weight_28_28;
wire signed[15:0]    spare_reg_psum_28_28;
wire signed[15:0]    spare_reg_weight_28_29;
wire signed[15:0]    spare_reg_psum_28_29;
wire signed[15:0]    spare_reg_weight_28_30;
wire signed[15:0]    spare_reg_psum_28_30;
wire signed[15:0]    spare_reg_weight_28_31;
wire signed[15:0]    spare_reg_psum_28_31;
wire signed[15:0]    spare_reg_weight_29_0;
wire signed[15:0]    spare_reg_psum_29_0;
wire signed[15:0]    spare_reg_weight_29_1;
wire signed[15:0]    spare_reg_psum_29_1;
wire signed[15:0]    spare_reg_weight_29_2;
wire signed[15:0]    spare_reg_psum_29_2;
wire signed[15:0]    spare_reg_weight_29_3;
wire signed[15:0]    spare_reg_psum_29_3;
wire signed[15:0]    spare_reg_weight_29_4;
wire signed[15:0]    spare_reg_psum_29_4;
wire signed[15:0]    spare_reg_weight_29_5;
wire signed[15:0]    spare_reg_psum_29_5;
wire signed[15:0]    spare_reg_weight_29_6;
wire signed[15:0]    spare_reg_psum_29_6;
wire signed[15:0]    spare_reg_weight_29_7;
wire signed[15:0]    spare_reg_psum_29_7;
wire signed[15:0]    spare_reg_weight_29_8;
wire signed[15:0]    spare_reg_psum_29_8;
wire signed[15:0]    spare_reg_weight_29_9;
wire signed[15:0]    spare_reg_psum_29_9;
wire signed[15:0]    spare_reg_weight_29_10;
wire signed[15:0]    spare_reg_psum_29_10;
wire signed[15:0]    spare_reg_weight_29_11;
wire signed[15:0]    spare_reg_psum_29_11;
wire signed[15:0]    spare_reg_weight_29_12;
wire signed[15:0]    spare_reg_psum_29_12;
wire signed[15:0]    spare_reg_weight_29_13;
wire signed[15:0]    spare_reg_psum_29_13;
wire signed[15:0]    spare_reg_weight_29_14;
wire signed[15:0]    spare_reg_psum_29_14;
wire signed[15:0]    spare_reg_weight_29_15;
wire signed[15:0]    spare_reg_psum_29_15;
wire signed[15:0]    spare_reg_weight_29_16;
wire signed[15:0]    spare_reg_psum_29_16;
wire signed[15:0]    spare_reg_weight_29_17;
wire signed[15:0]    spare_reg_psum_29_17;
wire signed[15:0]    spare_reg_weight_29_18;
wire signed[15:0]    spare_reg_psum_29_18;
wire signed[15:0]    spare_reg_weight_29_19;
wire signed[15:0]    spare_reg_psum_29_19;
wire signed[15:0]    spare_reg_weight_29_20;
wire signed[15:0]    spare_reg_psum_29_20;
wire signed[15:0]    spare_reg_weight_29_21;
wire signed[15:0]    spare_reg_psum_29_21;
wire signed[15:0]    spare_reg_weight_29_22;
wire signed[15:0]    spare_reg_psum_29_22;
wire signed[15:0]    spare_reg_weight_29_23;
wire signed[15:0]    spare_reg_psum_29_23;
wire signed[15:0]    spare_reg_weight_29_24;
wire signed[15:0]    spare_reg_psum_29_24;
wire signed[15:0]    spare_reg_weight_29_25;
wire signed[15:0]    spare_reg_psum_29_25;
wire signed[15:0]    spare_reg_weight_29_26;
wire signed[15:0]    spare_reg_psum_29_26;
wire signed[15:0]    spare_reg_weight_29_27;
wire signed[15:0]    spare_reg_psum_29_27;
wire signed[15:0]    spare_reg_weight_29_28;
wire signed[15:0]    spare_reg_psum_29_28;
wire signed[15:0]    spare_reg_weight_29_29;
wire signed[15:0]    spare_reg_psum_29_29;
wire signed[15:0]    spare_reg_weight_29_30;
wire signed[15:0]    spare_reg_psum_29_30;
wire signed[15:0]    spare_reg_weight_29_31;
wire signed[15:0]    spare_reg_psum_29_31;
wire signed[15:0]    spare_reg_weight_30_0;
wire signed[15:0]    spare_reg_psum_30_0;
wire signed[15:0]    spare_reg_weight_30_1;
wire signed[15:0]    spare_reg_psum_30_1;
wire signed[15:0]    spare_reg_weight_30_2;
wire signed[15:0]    spare_reg_psum_30_2;
wire signed[15:0]    spare_reg_weight_30_3;
wire signed[15:0]    spare_reg_psum_30_3;
wire signed[15:0]    spare_reg_weight_30_4;
wire signed[15:0]    spare_reg_psum_30_4;
wire signed[15:0]    spare_reg_weight_30_5;
wire signed[15:0]    spare_reg_psum_30_5;
wire signed[15:0]    spare_reg_weight_30_6;
wire signed[15:0]    spare_reg_psum_30_6;
wire signed[15:0]    spare_reg_weight_30_7;
wire signed[15:0]    spare_reg_psum_30_7;
wire signed[15:0]    spare_reg_weight_30_8;
wire signed[15:0]    spare_reg_psum_30_8;
wire signed[15:0]    spare_reg_weight_30_9;
wire signed[15:0]    spare_reg_psum_30_9;
wire signed[15:0]    spare_reg_weight_30_10;
wire signed[15:0]    spare_reg_psum_30_10;
wire signed[15:0]    spare_reg_weight_30_11;
wire signed[15:0]    spare_reg_psum_30_11;
wire signed[15:0]    spare_reg_weight_30_12;
wire signed[15:0]    spare_reg_psum_30_12;
wire signed[15:0]    spare_reg_weight_30_13;
wire signed[15:0]    spare_reg_psum_30_13;
wire signed[15:0]    spare_reg_weight_30_14;
wire signed[15:0]    spare_reg_psum_30_14;
wire signed[15:0]    spare_reg_weight_30_15;
wire signed[15:0]    spare_reg_psum_30_15;
wire signed[15:0]    spare_reg_weight_30_16;
wire signed[15:0]    spare_reg_psum_30_16;
wire signed[15:0]    spare_reg_weight_30_17;
wire signed[15:0]    spare_reg_psum_30_17;
wire signed[15:0]    spare_reg_weight_30_18;
wire signed[15:0]    spare_reg_psum_30_18;
wire signed[15:0]    spare_reg_weight_30_19;
wire signed[15:0]    spare_reg_psum_30_19;
wire signed[15:0]    spare_reg_weight_30_20;
wire signed[15:0]    spare_reg_psum_30_20;
wire signed[15:0]    spare_reg_weight_30_21;
wire signed[15:0]    spare_reg_psum_30_21;
wire signed[15:0]    spare_reg_weight_30_22;
wire signed[15:0]    spare_reg_psum_30_22;
wire signed[15:0]    spare_reg_weight_30_23;
wire signed[15:0]    spare_reg_psum_30_23;
wire signed[15:0]    spare_reg_weight_30_24;
wire signed[15:0]    spare_reg_psum_30_24;
wire signed[15:0]    spare_reg_weight_30_25;
wire signed[15:0]    spare_reg_psum_30_25;
wire signed[15:0]    spare_reg_weight_30_26;
wire signed[15:0]    spare_reg_psum_30_26;
wire signed[15:0]    spare_reg_weight_30_27;
wire signed[15:0]    spare_reg_psum_30_27;
wire signed[15:0]    spare_reg_weight_30_28;
wire signed[15:0]    spare_reg_psum_30_28;
wire signed[15:0]    spare_reg_weight_30_29;
wire signed[15:0]    spare_reg_psum_30_29;
wire signed[15:0]    spare_reg_weight_30_30;
wire signed[15:0]    spare_reg_psum_30_30;
wire signed[15:0]    spare_reg_weight_30_31;
wire signed[15:0]    spare_reg_psum_30_31;
wire signed[15:0]    spare_reg_weight_31_0;
wire signed[15:0]    spare_reg_psum_31_0;
wire signed[15:0]    spare_reg_weight_31_1;
wire signed[15:0]    spare_reg_psum_31_1;
wire signed[15:0]    spare_reg_weight_31_2;
wire signed[15:0]    spare_reg_psum_31_2;
wire signed[15:0]    spare_reg_weight_31_3;
wire signed[15:0]    spare_reg_psum_31_3;
wire signed[15:0]    spare_reg_weight_31_4;
wire signed[15:0]    spare_reg_psum_31_4;
wire signed[15:0]    spare_reg_weight_31_5;
wire signed[15:0]    spare_reg_psum_31_5;
wire signed[15:0]    spare_reg_weight_31_6;
wire signed[15:0]    spare_reg_psum_31_6;
wire signed[15:0]    spare_reg_weight_31_7;
wire signed[15:0]    spare_reg_psum_31_7;
wire signed[15:0]    spare_reg_weight_31_8;
wire signed[15:0]    spare_reg_psum_31_8;
wire signed[15:0]    spare_reg_weight_31_9;
wire signed[15:0]    spare_reg_psum_31_9;
wire signed[15:0]    spare_reg_weight_31_10;
wire signed[15:0]    spare_reg_psum_31_10;
wire signed[15:0]    spare_reg_weight_31_11;
wire signed[15:0]    spare_reg_psum_31_11;
wire signed[15:0]    spare_reg_weight_31_12;
wire signed[15:0]    spare_reg_psum_31_12;
wire signed[15:0]    spare_reg_weight_31_13;
wire signed[15:0]    spare_reg_psum_31_13;
wire signed[15:0]    spare_reg_weight_31_14;
wire signed[15:0]    spare_reg_psum_31_14;
wire signed[15:0]    spare_reg_weight_31_15;
wire signed[15:0]    spare_reg_psum_31_15;
wire signed[15:0]    spare_reg_weight_31_16;
wire signed[15:0]    spare_reg_psum_31_16;
wire signed[15:0]    spare_reg_weight_31_17;
wire signed[15:0]    spare_reg_psum_31_17;
wire signed[15:0]    spare_reg_weight_31_18;
wire signed[15:0]    spare_reg_psum_31_18;
wire signed[15:0]    spare_reg_weight_31_19;
wire signed[15:0]    spare_reg_psum_31_19;
wire signed[15:0]    spare_reg_weight_31_20;
wire signed[15:0]    spare_reg_psum_31_20;
wire signed[15:0]    spare_reg_weight_31_21;
wire signed[15:0]    spare_reg_psum_31_21;
wire signed[15:0]    spare_reg_weight_31_22;
wire signed[15:0]    spare_reg_psum_31_22;
wire signed[15:0]    spare_reg_weight_31_23;
wire signed[15:0]    spare_reg_psum_31_23;
wire signed[15:0]    spare_reg_weight_31_24;
wire signed[15:0]    spare_reg_psum_31_24;
wire signed[15:0]    spare_reg_weight_31_25;
wire signed[15:0]    spare_reg_psum_31_25;
wire signed[15:0]    spare_reg_weight_31_26;
wire signed[15:0]    spare_reg_psum_31_26;
wire signed[15:0]    spare_reg_weight_31_27;
wire signed[15:0]    spare_reg_psum_31_27;
wire signed[15:0]    spare_reg_weight_31_28;
wire signed[15:0]    spare_reg_psum_31_28;
wire signed[15:0]    spare_reg_weight_31_29;
wire signed[15:0]    spare_reg_psum_31_29;
wire signed[15:0]    spare_reg_weight_31_30;
wire signed[15:0]    spare_reg_psum_31_30;
wire signed[15:0]    spare_reg_weight_31_31;
wire signed[15:0]    spare_reg_psum_31_31;
output signed[15:0]   spare_out_psum_0;
output signed[15:0]   spare_out_psum_1;
output signed[15:0]   spare_out_psum_2;
output signed[15:0]   spare_out_psum_3;
output signed[15:0]   spare_out_psum_4;
output signed[15:0]   spare_out_psum_5;
output signed[15:0]   spare_out_psum_6;
output signed[15:0]   spare_out_psum_7;
output signed[15:0]   spare_out_psum_8;
output signed[15:0]   spare_out_psum_9;
output signed[15:0]   spare_out_psum_10;
output signed[15:0]   spare_out_psum_11;
output signed[15:0]   spare_out_psum_12;
output signed[15:0]   spare_out_psum_13;
output signed[15:0]   spare_out_psum_14;
output signed[15:0]   spare_out_psum_15;
output signed[15:0]   spare_out_psum_16;
output signed[15:0]   spare_out_psum_17;
output signed[15:0]   spare_out_psum_18;
output signed[15:0]   spare_out_psum_19;
output signed[15:0]   spare_out_psum_20;
output signed[15:0]   spare_out_psum_21;
output signed[15:0]   spare_out_psum_22;
output signed[15:0]   spare_out_psum_23;
output signed[15:0]   spare_out_psum_24;
output signed[15:0]   spare_out_psum_25;
output signed[15:0]   spare_out_psum_26;
output signed[15:0]   spare_out_psum_27;
output signed[15:0]   spare_out_psum_28;
output signed[15:0]   spare_out_psum_29;
output signed[15:0]   spare_out_psum_30;
output signed[15:0]   spare_out_psum_31;
assign spare_out_psum_0 =  spare_reg_psum_31_0;
assign spare_out_psum_1 =  spare_reg_psum_31_1;
assign spare_out_psum_2 =  spare_reg_psum_31_2;
assign spare_out_psum_3 =  spare_reg_psum_31_3;
assign spare_out_psum_4 =  spare_reg_psum_31_4;
assign spare_out_psum_5 =  spare_reg_psum_31_5;
assign spare_out_psum_6 =  spare_reg_psum_31_6;
assign spare_out_psum_7 =  spare_reg_psum_31_7;
assign spare_out_psum_8 =  spare_reg_psum_31_8;
assign spare_out_psum_9 =  spare_reg_psum_31_9;
assign spare_out_psum_10 =  spare_reg_psum_31_10;
assign spare_out_psum_11 =  spare_reg_psum_31_11;
assign spare_out_psum_12 =  spare_reg_psum_31_12;
assign spare_out_psum_13 =  spare_reg_psum_31_13;
assign spare_out_psum_14 =  spare_reg_psum_31_14;
assign spare_out_psum_15 =  spare_reg_psum_31_15;
assign spare_out_psum_16 =  spare_reg_psum_31_16;
assign spare_out_psum_17 =  spare_reg_psum_31_17;
assign spare_out_psum_18 =  spare_reg_psum_31_18;
assign spare_out_psum_19 =  spare_reg_psum_31_19;
assign spare_out_psum_20 =  spare_reg_psum_31_20;
assign spare_out_psum_21 =  spare_reg_psum_31_21;
assign spare_out_psum_22 =  spare_reg_psum_31_22;
assign spare_out_psum_23 =  spare_reg_psum_31_23;
assign spare_out_psum_24 =  spare_reg_psum_31_24;
assign spare_out_psum_25 =  spare_reg_psum_31_25;
assign spare_out_psum_26 =  spare_reg_psum_31_26;
assign spare_out_psum_27 =  spare_reg_psum_31_27;
assign spare_out_psum_28 =  spare_reg_psum_31_28;
assign spare_out_psum_29 =  spare_reg_psum_31_29;
assign spare_out_psum_30 =  spare_reg_psum_31_30;
assign spare_out_psum_31 =  spare_reg_psum_31_31;
PE X0_0( .activation_in(in_activation_0), .weight_in(in_weight_0), .partial_sum_in(in_psum_0), .reg_activation(spare_reg_activation_0_0), .reg_weight(spare_reg_weight_0_0), .reg_partial_sum(spare_reg_psum_0_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_1( .activation_in(spare_reg_activation_0_0), .weight_in(in_weight_1), .partial_sum_in(in_psum_1), .reg_activation(spare_reg_activation_0_1), .reg_weight(spare_reg_weight_0_1), .reg_partial_sum(spare_reg_psum_0_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_2( .activation_in(spare_reg_activation_0_1), .weight_in(in_weight_2), .partial_sum_in(in_psum_2), .reg_activation(spare_reg_activation_0_2), .reg_weight(spare_reg_weight_0_2), .reg_partial_sum(spare_reg_psum_0_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_3( .activation_in(spare_reg_activation_0_2), .weight_in(in_weight_3), .partial_sum_in(in_psum_3), .reg_activation(spare_reg_activation_0_3), .reg_weight(spare_reg_weight_0_3), .reg_partial_sum(spare_reg_psum_0_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_4( .activation_in(spare_reg_activation_0_3), .weight_in(in_weight_4), .partial_sum_in(in_psum_4), .reg_activation(spare_reg_activation_0_4), .reg_weight(spare_reg_weight_0_4), .reg_partial_sum(spare_reg_psum_0_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_5( .activation_in(spare_reg_activation_0_4), .weight_in(in_weight_5), .partial_sum_in(in_psum_5), .reg_activation(spare_reg_activation_0_5), .reg_weight(spare_reg_weight_0_5), .reg_partial_sum(spare_reg_psum_0_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_6( .activation_in(spare_reg_activation_0_5), .weight_in(in_weight_6), .partial_sum_in(in_psum_6), .reg_activation(spare_reg_activation_0_6), .reg_weight(spare_reg_weight_0_6), .reg_partial_sum(spare_reg_psum_0_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_7( .activation_in(spare_reg_activation_0_6), .weight_in(in_weight_7), .partial_sum_in(in_psum_7), .reg_activation(spare_reg_activation_0_7), .reg_weight(spare_reg_weight_0_7), .reg_partial_sum(spare_reg_psum_0_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_8( .activation_in(spare_reg_activation_0_7), .weight_in(in_weight_8), .partial_sum_in(in_psum_8), .reg_activation(spare_reg_activation_0_8), .reg_weight(spare_reg_weight_0_8), .reg_partial_sum(spare_reg_psum_0_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_9( .activation_in(spare_reg_activation_0_8), .weight_in(in_weight_9), .partial_sum_in(in_psum_9), .reg_activation(spare_reg_activation_0_9), .reg_weight(spare_reg_weight_0_9), .reg_partial_sum(spare_reg_psum_0_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_10( .activation_in(spare_reg_activation_0_9), .weight_in(in_weight_10), .partial_sum_in(in_psum_10), .reg_activation(spare_reg_activation_0_10), .reg_weight(spare_reg_weight_0_10), .reg_partial_sum(spare_reg_psum_0_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_11( .activation_in(spare_reg_activation_0_10), .weight_in(in_weight_11), .partial_sum_in(in_psum_11), .reg_activation(spare_reg_activation_0_11), .reg_weight(spare_reg_weight_0_11), .reg_partial_sum(spare_reg_psum_0_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_12( .activation_in(spare_reg_activation_0_11), .weight_in(in_weight_12), .partial_sum_in(in_psum_12), .reg_activation(spare_reg_activation_0_12), .reg_weight(spare_reg_weight_0_12), .reg_partial_sum(spare_reg_psum_0_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_13( .activation_in(spare_reg_activation_0_12), .weight_in(in_weight_13), .partial_sum_in(in_psum_13), .reg_activation(spare_reg_activation_0_13), .reg_weight(spare_reg_weight_0_13), .reg_partial_sum(spare_reg_psum_0_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_14( .activation_in(spare_reg_activation_0_13), .weight_in(in_weight_14), .partial_sum_in(in_psum_14), .reg_activation(spare_reg_activation_0_14), .reg_weight(spare_reg_weight_0_14), .reg_partial_sum(spare_reg_psum_0_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_15( .activation_in(spare_reg_activation_0_14), .weight_in(in_weight_15), .partial_sum_in(in_psum_15), .reg_activation(spare_reg_activation_0_15), .reg_weight(spare_reg_weight_0_15), .reg_partial_sum(spare_reg_psum_0_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_16( .activation_in(spare_reg_activation_0_15), .weight_in(in_weight_16), .partial_sum_in(in_psum_16), .reg_activation(spare_reg_activation_0_16), .reg_weight(spare_reg_weight_0_16), .reg_partial_sum(spare_reg_psum_0_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_17( .activation_in(spare_reg_activation_0_16), .weight_in(in_weight_17), .partial_sum_in(in_psum_17), .reg_activation(spare_reg_activation_0_17), .reg_weight(spare_reg_weight_0_17), .reg_partial_sum(spare_reg_psum_0_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_18( .activation_in(spare_reg_activation_0_17), .weight_in(in_weight_18), .partial_sum_in(in_psum_18), .reg_activation(spare_reg_activation_0_18), .reg_weight(spare_reg_weight_0_18), .reg_partial_sum(spare_reg_psum_0_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_19( .activation_in(spare_reg_activation_0_18), .weight_in(in_weight_19), .partial_sum_in(in_psum_19), .reg_activation(spare_reg_activation_0_19), .reg_weight(spare_reg_weight_0_19), .reg_partial_sum(spare_reg_psum_0_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_20( .activation_in(spare_reg_activation_0_19), .weight_in(in_weight_20), .partial_sum_in(in_psum_20), .reg_activation(spare_reg_activation_0_20), .reg_weight(spare_reg_weight_0_20), .reg_partial_sum(spare_reg_psum_0_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_21( .activation_in(spare_reg_activation_0_20), .weight_in(in_weight_21), .partial_sum_in(in_psum_21), .reg_activation(spare_reg_activation_0_21), .reg_weight(spare_reg_weight_0_21), .reg_partial_sum(spare_reg_psum_0_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_22( .activation_in(spare_reg_activation_0_21), .weight_in(in_weight_22), .partial_sum_in(in_psum_22), .reg_activation(spare_reg_activation_0_22), .reg_weight(spare_reg_weight_0_22), .reg_partial_sum(spare_reg_psum_0_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_23( .activation_in(spare_reg_activation_0_22), .weight_in(in_weight_23), .partial_sum_in(in_psum_23), .reg_activation(spare_reg_activation_0_23), .reg_weight(spare_reg_weight_0_23), .reg_partial_sum(spare_reg_psum_0_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_24( .activation_in(spare_reg_activation_0_23), .weight_in(in_weight_24), .partial_sum_in(in_psum_24), .reg_activation(spare_reg_activation_0_24), .reg_weight(spare_reg_weight_0_24), .reg_partial_sum(spare_reg_psum_0_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_25( .activation_in(spare_reg_activation_0_24), .weight_in(in_weight_25), .partial_sum_in(in_psum_25), .reg_activation(spare_reg_activation_0_25), .reg_weight(spare_reg_weight_0_25), .reg_partial_sum(spare_reg_psum_0_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_26( .activation_in(spare_reg_activation_0_25), .weight_in(in_weight_26), .partial_sum_in(in_psum_26), .reg_activation(spare_reg_activation_0_26), .reg_weight(spare_reg_weight_0_26), .reg_partial_sum(spare_reg_psum_0_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_27( .activation_in(spare_reg_activation_0_26), .weight_in(in_weight_27), .partial_sum_in(in_psum_27), .reg_activation(spare_reg_activation_0_27), .reg_weight(spare_reg_weight_0_27), .reg_partial_sum(spare_reg_psum_0_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_28( .activation_in(spare_reg_activation_0_27), .weight_in(in_weight_28), .partial_sum_in(in_psum_28), .reg_activation(spare_reg_activation_0_28), .reg_weight(spare_reg_weight_0_28), .reg_partial_sum(spare_reg_psum_0_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_29( .activation_in(spare_reg_activation_0_28), .weight_in(in_weight_29), .partial_sum_in(in_psum_29), .reg_activation(spare_reg_activation_0_29), .reg_weight(spare_reg_weight_0_29), .reg_partial_sum(spare_reg_psum_0_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_30( .activation_in(spare_reg_activation_0_29), .weight_in(in_weight_30), .partial_sum_in(in_psum_30), .reg_activation(spare_reg_activation_0_30), .reg_weight(spare_reg_weight_0_30), .reg_partial_sum(spare_reg_psum_0_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X0_31( .activation_in(spare_reg_activation_0_30), .weight_in(in_weight_31), .partial_sum_in(in_psum_31), .reg_weight(spare_reg_weight_0_31), .reg_partial_sum(spare_reg_psum_0_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_0( .activation_in(in_activation_1), .weight_in(spare_reg_weight_0_0), .partial_sum_in(spare_reg_psum_0_0), .reg_activation(spare_reg_activation_1_0), .reg_weight(spare_reg_weight_1_0), .reg_partial_sum(spare_reg_psum_1_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_1( .activation_in(spare_reg_activation_1_0), .weight_in(spare_reg_weight_0_1), .partial_sum_in(spare_reg_psum_0_1), .reg_activation(spare_reg_activation_1_1), .reg_weight(spare_reg_weight_1_1), .reg_partial_sum(spare_reg_psum_1_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_2( .activation_in(spare_reg_activation_1_1), .weight_in(spare_reg_weight_0_2), .partial_sum_in(spare_reg_psum_0_2), .reg_activation(spare_reg_activation_1_2), .reg_weight(spare_reg_weight_1_2), .reg_partial_sum(spare_reg_psum_1_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_3( .activation_in(spare_reg_activation_1_2), .weight_in(spare_reg_weight_0_3), .partial_sum_in(spare_reg_psum_0_3), .reg_activation(spare_reg_activation_1_3), .reg_weight(spare_reg_weight_1_3), .reg_partial_sum(spare_reg_psum_1_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_4( .activation_in(spare_reg_activation_1_3), .weight_in(spare_reg_weight_0_4), .partial_sum_in(spare_reg_psum_0_4), .reg_activation(spare_reg_activation_1_4), .reg_weight(spare_reg_weight_1_4), .reg_partial_sum(spare_reg_psum_1_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_5( .activation_in(spare_reg_activation_1_4), .weight_in(spare_reg_weight_0_5), .partial_sum_in(spare_reg_psum_0_5), .reg_activation(spare_reg_activation_1_5), .reg_weight(spare_reg_weight_1_5), .reg_partial_sum(spare_reg_psum_1_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_6( .activation_in(spare_reg_activation_1_5), .weight_in(spare_reg_weight_0_6), .partial_sum_in(spare_reg_psum_0_6), .reg_activation(spare_reg_activation_1_6), .reg_weight(spare_reg_weight_1_6), .reg_partial_sum(spare_reg_psum_1_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_7( .activation_in(spare_reg_activation_1_6), .weight_in(spare_reg_weight_0_7), .partial_sum_in(spare_reg_psum_0_7), .reg_activation(spare_reg_activation_1_7), .reg_weight(spare_reg_weight_1_7), .reg_partial_sum(spare_reg_psum_1_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_8( .activation_in(spare_reg_activation_1_7), .weight_in(spare_reg_weight_0_8), .partial_sum_in(spare_reg_psum_0_8), .reg_activation(spare_reg_activation_1_8), .reg_weight(spare_reg_weight_1_8), .reg_partial_sum(spare_reg_psum_1_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_9( .activation_in(spare_reg_activation_1_8), .weight_in(spare_reg_weight_0_9), .partial_sum_in(spare_reg_psum_0_9), .reg_activation(spare_reg_activation_1_9), .reg_weight(spare_reg_weight_1_9), .reg_partial_sum(spare_reg_psum_1_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_10( .activation_in(spare_reg_activation_1_9), .weight_in(spare_reg_weight_0_10), .partial_sum_in(spare_reg_psum_0_10), .reg_activation(spare_reg_activation_1_10), .reg_weight(spare_reg_weight_1_10), .reg_partial_sum(spare_reg_psum_1_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_11( .activation_in(spare_reg_activation_1_10), .weight_in(spare_reg_weight_0_11), .partial_sum_in(spare_reg_psum_0_11), .reg_activation(spare_reg_activation_1_11), .reg_weight(spare_reg_weight_1_11), .reg_partial_sum(spare_reg_psum_1_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_12( .activation_in(spare_reg_activation_1_11), .weight_in(spare_reg_weight_0_12), .partial_sum_in(spare_reg_psum_0_12), .reg_activation(spare_reg_activation_1_12), .reg_weight(spare_reg_weight_1_12), .reg_partial_sum(spare_reg_psum_1_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_13( .activation_in(spare_reg_activation_1_12), .weight_in(spare_reg_weight_0_13), .partial_sum_in(spare_reg_psum_0_13), .reg_activation(spare_reg_activation_1_13), .reg_weight(spare_reg_weight_1_13), .reg_partial_sum(spare_reg_psum_1_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_14( .activation_in(spare_reg_activation_1_13), .weight_in(spare_reg_weight_0_14), .partial_sum_in(spare_reg_psum_0_14), .reg_activation(spare_reg_activation_1_14), .reg_weight(spare_reg_weight_1_14), .reg_partial_sum(spare_reg_psum_1_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_15( .activation_in(spare_reg_activation_1_14), .weight_in(spare_reg_weight_0_15), .partial_sum_in(spare_reg_psum_0_15), .reg_activation(spare_reg_activation_1_15), .reg_weight(spare_reg_weight_1_15), .reg_partial_sum(spare_reg_psum_1_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_16( .activation_in(spare_reg_activation_1_15), .weight_in(spare_reg_weight_0_16), .partial_sum_in(spare_reg_psum_0_16), .reg_activation(spare_reg_activation_1_16), .reg_weight(spare_reg_weight_1_16), .reg_partial_sum(spare_reg_psum_1_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_17( .activation_in(spare_reg_activation_1_16), .weight_in(spare_reg_weight_0_17), .partial_sum_in(spare_reg_psum_0_17), .reg_activation(spare_reg_activation_1_17), .reg_weight(spare_reg_weight_1_17), .reg_partial_sum(spare_reg_psum_1_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_18( .activation_in(spare_reg_activation_1_17), .weight_in(spare_reg_weight_0_18), .partial_sum_in(spare_reg_psum_0_18), .reg_activation(spare_reg_activation_1_18), .reg_weight(spare_reg_weight_1_18), .reg_partial_sum(spare_reg_psum_1_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_19( .activation_in(spare_reg_activation_1_18), .weight_in(spare_reg_weight_0_19), .partial_sum_in(spare_reg_psum_0_19), .reg_activation(spare_reg_activation_1_19), .reg_weight(spare_reg_weight_1_19), .reg_partial_sum(spare_reg_psum_1_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_20( .activation_in(spare_reg_activation_1_19), .weight_in(spare_reg_weight_0_20), .partial_sum_in(spare_reg_psum_0_20), .reg_activation(spare_reg_activation_1_20), .reg_weight(spare_reg_weight_1_20), .reg_partial_sum(spare_reg_psum_1_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_21( .activation_in(spare_reg_activation_1_20), .weight_in(spare_reg_weight_0_21), .partial_sum_in(spare_reg_psum_0_21), .reg_activation(spare_reg_activation_1_21), .reg_weight(spare_reg_weight_1_21), .reg_partial_sum(spare_reg_psum_1_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_22( .activation_in(spare_reg_activation_1_21), .weight_in(spare_reg_weight_0_22), .partial_sum_in(spare_reg_psum_0_22), .reg_activation(spare_reg_activation_1_22), .reg_weight(spare_reg_weight_1_22), .reg_partial_sum(spare_reg_psum_1_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_23( .activation_in(spare_reg_activation_1_22), .weight_in(spare_reg_weight_0_23), .partial_sum_in(spare_reg_psum_0_23), .reg_activation(spare_reg_activation_1_23), .reg_weight(spare_reg_weight_1_23), .reg_partial_sum(spare_reg_psum_1_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_24( .activation_in(spare_reg_activation_1_23), .weight_in(spare_reg_weight_0_24), .partial_sum_in(spare_reg_psum_0_24), .reg_activation(spare_reg_activation_1_24), .reg_weight(spare_reg_weight_1_24), .reg_partial_sum(spare_reg_psum_1_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_25( .activation_in(spare_reg_activation_1_24), .weight_in(spare_reg_weight_0_25), .partial_sum_in(spare_reg_psum_0_25), .reg_activation(spare_reg_activation_1_25), .reg_weight(spare_reg_weight_1_25), .reg_partial_sum(spare_reg_psum_1_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_26( .activation_in(spare_reg_activation_1_25), .weight_in(spare_reg_weight_0_26), .partial_sum_in(spare_reg_psum_0_26), .reg_activation(spare_reg_activation_1_26), .reg_weight(spare_reg_weight_1_26), .reg_partial_sum(spare_reg_psum_1_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_27( .activation_in(spare_reg_activation_1_26), .weight_in(spare_reg_weight_0_27), .partial_sum_in(spare_reg_psum_0_27), .reg_activation(spare_reg_activation_1_27), .reg_weight(spare_reg_weight_1_27), .reg_partial_sum(spare_reg_psum_1_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_28( .activation_in(spare_reg_activation_1_27), .weight_in(spare_reg_weight_0_28), .partial_sum_in(spare_reg_psum_0_28), .reg_activation(spare_reg_activation_1_28), .reg_weight(spare_reg_weight_1_28), .reg_partial_sum(spare_reg_psum_1_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_29( .activation_in(spare_reg_activation_1_28), .weight_in(spare_reg_weight_0_29), .partial_sum_in(spare_reg_psum_0_29), .reg_activation(spare_reg_activation_1_29), .reg_weight(spare_reg_weight_1_29), .reg_partial_sum(spare_reg_psum_1_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_30( .activation_in(spare_reg_activation_1_29), .weight_in(spare_reg_weight_0_30), .partial_sum_in(spare_reg_psum_0_30), .reg_activation(spare_reg_activation_1_30), .reg_weight(spare_reg_weight_1_30), .reg_partial_sum(spare_reg_psum_1_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X1_31( .activation_in(spare_reg_activation_1_30), .weight_in(spare_reg_weight_0_31), .partial_sum_in(spare_reg_psum_0_31), .reg_weight(spare_reg_weight_1_31), .reg_partial_sum(spare_reg_psum_1_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_0( .activation_in(in_activation_2), .weight_in(spare_reg_weight_1_0), .partial_sum_in(spare_reg_psum_1_0), .reg_activation(spare_reg_activation_2_0), .reg_weight(spare_reg_weight_2_0), .reg_partial_sum(spare_reg_psum_2_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_1( .activation_in(spare_reg_activation_2_0), .weight_in(spare_reg_weight_1_1), .partial_sum_in(spare_reg_psum_1_1), .reg_activation(spare_reg_activation_2_1), .reg_weight(spare_reg_weight_2_1), .reg_partial_sum(spare_reg_psum_2_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_2( .activation_in(spare_reg_activation_2_1), .weight_in(spare_reg_weight_1_2), .partial_sum_in(spare_reg_psum_1_2), .reg_activation(spare_reg_activation_2_2), .reg_weight(spare_reg_weight_2_2), .reg_partial_sum(spare_reg_psum_2_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_3( .activation_in(spare_reg_activation_2_2), .weight_in(spare_reg_weight_1_3), .partial_sum_in(spare_reg_psum_1_3), .reg_activation(spare_reg_activation_2_3), .reg_weight(spare_reg_weight_2_3), .reg_partial_sum(spare_reg_psum_2_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_4( .activation_in(spare_reg_activation_2_3), .weight_in(spare_reg_weight_1_4), .partial_sum_in(spare_reg_psum_1_4), .reg_activation(spare_reg_activation_2_4), .reg_weight(spare_reg_weight_2_4), .reg_partial_sum(spare_reg_psum_2_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_5( .activation_in(spare_reg_activation_2_4), .weight_in(spare_reg_weight_1_5), .partial_sum_in(spare_reg_psum_1_5), .reg_activation(spare_reg_activation_2_5), .reg_weight(spare_reg_weight_2_5), .reg_partial_sum(spare_reg_psum_2_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_6( .activation_in(spare_reg_activation_2_5), .weight_in(spare_reg_weight_1_6), .partial_sum_in(spare_reg_psum_1_6), .reg_activation(spare_reg_activation_2_6), .reg_weight(spare_reg_weight_2_6), .reg_partial_sum(spare_reg_psum_2_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_7( .activation_in(spare_reg_activation_2_6), .weight_in(spare_reg_weight_1_7), .partial_sum_in(spare_reg_psum_1_7), .reg_activation(spare_reg_activation_2_7), .reg_weight(spare_reg_weight_2_7), .reg_partial_sum(spare_reg_psum_2_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_8( .activation_in(spare_reg_activation_2_7), .weight_in(spare_reg_weight_1_8), .partial_sum_in(spare_reg_psum_1_8), .reg_activation(spare_reg_activation_2_8), .reg_weight(spare_reg_weight_2_8), .reg_partial_sum(spare_reg_psum_2_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_9( .activation_in(spare_reg_activation_2_8), .weight_in(spare_reg_weight_1_9), .partial_sum_in(spare_reg_psum_1_9), .reg_activation(spare_reg_activation_2_9), .reg_weight(spare_reg_weight_2_9), .reg_partial_sum(spare_reg_psum_2_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_10( .activation_in(spare_reg_activation_2_9), .weight_in(spare_reg_weight_1_10), .partial_sum_in(spare_reg_psum_1_10), .reg_activation(spare_reg_activation_2_10), .reg_weight(spare_reg_weight_2_10), .reg_partial_sum(spare_reg_psum_2_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_11( .activation_in(spare_reg_activation_2_10), .weight_in(spare_reg_weight_1_11), .partial_sum_in(spare_reg_psum_1_11), .reg_activation(spare_reg_activation_2_11), .reg_weight(spare_reg_weight_2_11), .reg_partial_sum(spare_reg_psum_2_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_12( .activation_in(spare_reg_activation_2_11), .weight_in(spare_reg_weight_1_12), .partial_sum_in(spare_reg_psum_1_12), .reg_activation(spare_reg_activation_2_12), .reg_weight(spare_reg_weight_2_12), .reg_partial_sum(spare_reg_psum_2_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_13( .activation_in(spare_reg_activation_2_12), .weight_in(spare_reg_weight_1_13), .partial_sum_in(spare_reg_psum_1_13), .reg_activation(spare_reg_activation_2_13), .reg_weight(spare_reg_weight_2_13), .reg_partial_sum(spare_reg_psum_2_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_14( .activation_in(spare_reg_activation_2_13), .weight_in(spare_reg_weight_1_14), .partial_sum_in(spare_reg_psum_1_14), .reg_activation(spare_reg_activation_2_14), .reg_weight(spare_reg_weight_2_14), .reg_partial_sum(spare_reg_psum_2_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_15( .activation_in(spare_reg_activation_2_14), .weight_in(spare_reg_weight_1_15), .partial_sum_in(spare_reg_psum_1_15), .reg_activation(spare_reg_activation_2_15), .reg_weight(spare_reg_weight_2_15), .reg_partial_sum(spare_reg_psum_2_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_16( .activation_in(spare_reg_activation_2_15), .weight_in(spare_reg_weight_1_16), .partial_sum_in(spare_reg_psum_1_16), .reg_activation(spare_reg_activation_2_16), .reg_weight(spare_reg_weight_2_16), .reg_partial_sum(spare_reg_psum_2_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_17( .activation_in(spare_reg_activation_2_16), .weight_in(spare_reg_weight_1_17), .partial_sum_in(spare_reg_psum_1_17), .reg_activation(spare_reg_activation_2_17), .reg_weight(spare_reg_weight_2_17), .reg_partial_sum(spare_reg_psum_2_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_18( .activation_in(spare_reg_activation_2_17), .weight_in(spare_reg_weight_1_18), .partial_sum_in(spare_reg_psum_1_18), .reg_activation(spare_reg_activation_2_18), .reg_weight(spare_reg_weight_2_18), .reg_partial_sum(spare_reg_psum_2_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_19( .activation_in(spare_reg_activation_2_18), .weight_in(spare_reg_weight_1_19), .partial_sum_in(spare_reg_psum_1_19), .reg_activation(spare_reg_activation_2_19), .reg_weight(spare_reg_weight_2_19), .reg_partial_sum(spare_reg_psum_2_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_20( .activation_in(spare_reg_activation_2_19), .weight_in(spare_reg_weight_1_20), .partial_sum_in(spare_reg_psum_1_20), .reg_activation(spare_reg_activation_2_20), .reg_weight(spare_reg_weight_2_20), .reg_partial_sum(spare_reg_psum_2_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_21( .activation_in(spare_reg_activation_2_20), .weight_in(spare_reg_weight_1_21), .partial_sum_in(spare_reg_psum_1_21), .reg_activation(spare_reg_activation_2_21), .reg_weight(spare_reg_weight_2_21), .reg_partial_sum(spare_reg_psum_2_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_22( .activation_in(spare_reg_activation_2_21), .weight_in(spare_reg_weight_1_22), .partial_sum_in(spare_reg_psum_1_22), .reg_activation(spare_reg_activation_2_22), .reg_weight(spare_reg_weight_2_22), .reg_partial_sum(spare_reg_psum_2_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_23( .activation_in(spare_reg_activation_2_22), .weight_in(spare_reg_weight_1_23), .partial_sum_in(spare_reg_psum_1_23), .reg_activation(spare_reg_activation_2_23), .reg_weight(spare_reg_weight_2_23), .reg_partial_sum(spare_reg_psum_2_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_24( .activation_in(spare_reg_activation_2_23), .weight_in(spare_reg_weight_1_24), .partial_sum_in(spare_reg_psum_1_24), .reg_activation(spare_reg_activation_2_24), .reg_weight(spare_reg_weight_2_24), .reg_partial_sum(spare_reg_psum_2_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_25( .activation_in(spare_reg_activation_2_24), .weight_in(spare_reg_weight_1_25), .partial_sum_in(spare_reg_psum_1_25), .reg_activation(spare_reg_activation_2_25), .reg_weight(spare_reg_weight_2_25), .reg_partial_sum(spare_reg_psum_2_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_26( .activation_in(spare_reg_activation_2_25), .weight_in(spare_reg_weight_1_26), .partial_sum_in(spare_reg_psum_1_26), .reg_activation(spare_reg_activation_2_26), .reg_weight(spare_reg_weight_2_26), .reg_partial_sum(spare_reg_psum_2_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_27( .activation_in(spare_reg_activation_2_26), .weight_in(spare_reg_weight_1_27), .partial_sum_in(spare_reg_psum_1_27), .reg_activation(spare_reg_activation_2_27), .reg_weight(spare_reg_weight_2_27), .reg_partial_sum(spare_reg_psum_2_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_28( .activation_in(spare_reg_activation_2_27), .weight_in(spare_reg_weight_1_28), .partial_sum_in(spare_reg_psum_1_28), .reg_activation(spare_reg_activation_2_28), .reg_weight(spare_reg_weight_2_28), .reg_partial_sum(spare_reg_psum_2_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_29( .activation_in(spare_reg_activation_2_28), .weight_in(spare_reg_weight_1_29), .partial_sum_in(spare_reg_psum_1_29), .reg_activation(spare_reg_activation_2_29), .reg_weight(spare_reg_weight_2_29), .reg_partial_sum(spare_reg_psum_2_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_30( .activation_in(spare_reg_activation_2_29), .weight_in(spare_reg_weight_1_30), .partial_sum_in(spare_reg_psum_1_30), .reg_activation(spare_reg_activation_2_30), .reg_weight(spare_reg_weight_2_30), .reg_partial_sum(spare_reg_psum_2_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X2_31( .activation_in(spare_reg_activation_2_30), .weight_in(spare_reg_weight_1_31), .partial_sum_in(spare_reg_psum_1_31), .reg_weight(spare_reg_weight_2_31), .reg_partial_sum(spare_reg_psum_2_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_0( .activation_in(in_activation_3), .weight_in(spare_reg_weight_2_0), .partial_sum_in(spare_reg_psum_2_0), .reg_activation(spare_reg_activation_3_0), .reg_weight(spare_reg_weight_3_0), .reg_partial_sum(spare_reg_psum_3_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_1( .activation_in(spare_reg_activation_3_0), .weight_in(spare_reg_weight_2_1), .partial_sum_in(spare_reg_psum_2_1), .reg_activation(spare_reg_activation_3_1), .reg_weight(spare_reg_weight_3_1), .reg_partial_sum(spare_reg_psum_3_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_2( .activation_in(spare_reg_activation_3_1), .weight_in(spare_reg_weight_2_2), .partial_sum_in(spare_reg_psum_2_2), .reg_activation(spare_reg_activation_3_2), .reg_weight(spare_reg_weight_3_2), .reg_partial_sum(spare_reg_psum_3_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_3( .activation_in(spare_reg_activation_3_2), .weight_in(spare_reg_weight_2_3), .partial_sum_in(spare_reg_psum_2_3), .reg_activation(spare_reg_activation_3_3), .reg_weight(spare_reg_weight_3_3), .reg_partial_sum(spare_reg_psum_3_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_4( .activation_in(spare_reg_activation_3_3), .weight_in(spare_reg_weight_2_4), .partial_sum_in(spare_reg_psum_2_4), .reg_activation(spare_reg_activation_3_4), .reg_weight(spare_reg_weight_3_4), .reg_partial_sum(spare_reg_psum_3_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_5( .activation_in(spare_reg_activation_3_4), .weight_in(spare_reg_weight_2_5), .partial_sum_in(spare_reg_psum_2_5), .reg_activation(spare_reg_activation_3_5), .reg_weight(spare_reg_weight_3_5), .reg_partial_sum(spare_reg_psum_3_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_6( .activation_in(spare_reg_activation_3_5), .weight_in(spare_reg_weight_2_6), .partial_sum_in(spare_reg_psum_2_6), .reg_activation(spare_reg_activation_3_6), .reg_weight(spare_reg_weight_3_6), .reg_partial_sum(spare_reg_psum_3_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_7( .activation_in(spare_reg_activation_3_6), .weight_in(spare_reg_weight_2_7), .partial_sum_in(spare_reg_psum_2_7), .reg_activation(spare_reg_activation_3_7), .reg_weight(spare_reg_weight_3_7), .reg_partial_sum(spare_reg_psum_3_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_8( .activation_in(spare_reg_activation_3_7), .weight_in(spare_reg_weight_2_8), .partial_sum_in(spare_reg_psum_2_8), .reg_activation(spare_reg_activation_3_8), .reg_weight(spare_reg_weight_3_8), .reg_partial_sum(spare_reg_psum_3_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_9( .activation_in(spare_reg_activation_3_8), .weight_in(spare_reg_weight_2_9), .partial_sum_in(spare_reg_psum_2_9), .reg_activation(spare_reg_activation_3_9), .reg_weight(spare_reg_weight_3_9), .reg_partial_sum(spare_reg_psum_3_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_10( .activation_in(spare_reg_activation_3_9), .weight_in(spare_reg_weight_2_10), .partial_sum_in(spare_reg_psum_2_10), .reg_activation(spare_reg_activation_3_10), .reg_weight(spare_reg_weight_3_10), .reg_partial_sum(spare_reg_psum_3_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_11( .activation_in(spare_reg_activation_3_10), .weight_in(spare_reg_weight_2_11), .partial_sum_in(spare_reg_psum_2_11), .reg_activation(spare_reg_activation_3_11), .reg_weight(spare_reg_weight_3_11), .reg_partial_sum(spare_reg_psum_3_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_12( .activation_in(spare_reg_activation_3_11), .weight_in(spare_reg_weight_2_12), .partial_sum_in(spare_reg_psum_2_12), .reg_activation(spare_reg_activation_3_12), .reg_weight(spare_reg_weight_3_12), .reg_partial_sum(spare_reg_psum_3_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_13( .activation_in(spare_reg_activation_3_12), .weight_in(spare_reg_weight_2_13), .partial_sum_in(spare_reg_psum_2_13), .reg_activation(spare_reg_activation_3_13), .reg_weight(spare_reg_weight_3_13), .reg_partial_sum(spare_reg_psum_3_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_14( .activation_in(spare_reg_activation_3_13), .weight_in(spare_reg_weight_2_14), .partial_sum_in(spare_reg_psum_2_14), .reg_activation(spare_reg_activation_3_14), .reg_weight(spare_reg_weight_3_14), .reg_partial_sum(spare_reg_psum_3_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_15( .activation_in(spare_reg_activation_3_14), .weight_in(spare_reg_weight_2_15), .partial_sum_in(spare_reg_psum_2_15), .reg_activation(spare_reg_activation_3_15), .reg_weight(spare_reg_weight_3_15), .reg_partial_sum(spare_reg_psum_3_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_16( .activation_in(spare_reg_activation_3_15), .weight_in(spare_reg_weight_2_16), .partial_sum_in(spare_reg_psum_2_16), .reg_activation(spare_reg_activation_3_16), .reg_weight(spare_reg_weight_3_16), .reg_partial_sum(spare_reg_psum_3_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_17( .activation_in(spare_reg_activation_3_16), .weight_in(spare_reg_weight_2_17), .partial_sum_in(spare_reg_psum_2_17), .reg_activation(spare_reg_activation_3_17), .reg_weight(spare_reg_weight_3_17), .reg_partial_sum(spare_reg_psum_3_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_18( .activation_in(spare_reg_activation_3_17), .weight_in(spare_reg_weight_2_18), .partial_sum_in(spare_reg_psum_2_18), .reg_activation(spare_reg_activation_3_18), .reg_weight(spare_reg_weight_3_18), .reg_partial_sum(spare_reg_psum_3_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_19( .activation_in(spare_reg_activation_3_18), .weight_in(spare_reg_weight_2_19), .partial_sum_in(spare_reg_psum_2_19), .reg_activation(spare_reg_activation_3_19), .reg_weight(spare_reg_weight_3_19), .reg_partial_sum(spare_reg_psum_3_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_20( .activation_in(spare_reg_activation_3_19), .weight_in(spare_reg_weight_2_20), .partial_sum_in(spare_reg_psum_2_20), .reg_activation(spare_reg_activation_3_20), .reg_weight(spare_reg_weight_3_20), .reg_partial_sum(spare_reg_psum_3_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_21( .activation_in(spare_reg_activation_3_20), .weight_in(spare_reg_weight_2_21), .partial_sum_in(spare_reg_psum_2_21), .reg_activation(spare_reg_activation_3_21), .reg_weight(spare_reg_weight_3_21), .reg_partial_sum(spare_reg_psum_3_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_22( .activation_in(spare_reg_activation_3_21), .weight_in(spare_reg_weight_2_22), .partial_sum_in(spare_reg_psum_2_22), .reg_activation(spare_reg_activation_3_22), .reg_weight(spare_reg_weight_3_22), .reg_partial_sum(spare_reg_psum_3_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_23( .activation_in(spare_reg_activation_3_22), .weight_in(spare_reg_weight_2_23), .partial_sum_in(spare_reg_psum_2_23), .reg_activation(spare_reg_activation_3_23), .reg_weight(spare_reg_weight_3_23), .reg_partial_sum(spare_reg_psum_3_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_24( .activation_in(spare_reg_activation_3_23), .weight_in(spare_reg_weight_2_24), .partial_sum_in(spare_reg_psum_2_24), .reg_activation(spare_reg_activation_3_24), .reg_weight(spare_reg_weight_3_24), .reg_partial_sum(spare_reg_psum_3_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_25( .activation_in(spare_reg_activation_3_24), .weight_in(spare_reg_weight_2_25), .partial_sum_in(spare_reg_psum_2_25), .reg_activation(spare_reg_activation_3_25), .reg_weight(spare_reg_weight_3_25), .reg_partial_sum(spare_reg_psum_3_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_26( .activation_in(spare_reg_activation_3_25), .weight_in(spare_reg_weight_2_26), .partial_sum_in(spare_reg_psum_2_26), .reg_activation(spare_reg_activation_3_26), .reg_weight(spare_reg_weight_3_26), .reg_partial_sum(spare_reg_psum_3_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_27( .activation_in(spare_reg_activation_3_26), .weight_in(spare_reg_weight_2_27), .partial_sum_in(spare_reg_psum_2_27), .reg_activation(spare_reg_activation_3_27), .reg_weight(spare_reg_weight_3_27), .reg_partial_sum(spare_reg_psum_3_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_28( .activation_in(spare_reg_activation_3_27), .weight_in(spare_reg_weight_2_28), .partial_sum_in(spare_reg_psum_2_28), .reg_activation(spare_reg_activation_3_28), .reg_weight(spare_reg_weight_3_28), .reg_partial_sum(spare_reg_psum_3_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_29( .activation_in(spare_reg_activation_3_28), .weight_in(spare_reg_weight_2_29), .partial_sum_in(spare_reg_psum_2_29), .reg_activation(spare_reg_activation_3_29), .reg_weight(spare_reg_weight_3_29), .reg_partial_sum(spare_reg_psum_3_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_30( .activation_in(spare_reg_activation_3_29), .weight_in(spare_reg_weight_2_30), .partial_sum_in(spare_reg_psum_2_30), .reg_activation(spare_reg_activation_3_30), .reg_weight(spare_reg_weight_3_30), .reg_partial_sum(spare_reg_psum_3_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X3_31( .activation_in(spare_reg_activation_3_30), .weight_in(spare_reg_weight_2_31), .partial_sum_in(spare_reg_psum_2_31), .reg_weight(spare_reg_weight_3_31), .reg_partial_sum(spare_reg_psum_3_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_0( .activation_in(in_activation_4), .weight_in(spare_reg_weight_3_0), .partial_sum_in(spare_reg_psum_3_0), .reg_activation(spare_reg_activation_4_0), .reg_weight(spare_reg_weight_4_0), .reg_partial_sum(spare_reg_psum_4_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_1( .activation_in(spare_reg_activation_4_0), .weight_in(spare_reg_weight_3_1), .partial_sum_in(spare_reg_psum_3_1), .reg_activation(spare_reg_activation_4_1), .reg_weight(spare_reg_weight_4_1), .reg_partial_sum(spare_reg_psum_4_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_2( .activation_in(spare_reg_activation_4_1), .weight_in(spare_reg_weight_3_2), .partial_sum_in(spare_reg_psum_3_2), .reg_activation(spare_reg_activation_4_2), .reg_weight(spare_reg_weight_4_2), .reg_partial_sum(spare_reg_psum_4_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_3( .activation_in(spare_reg_activation_4_2), .weight_in(spare_reg_weight_3_3), .partial_sum_in(spare_reg_psum_3_3), .reg_activation(spare_reg_activation_4_3), .reg_weight(spare_reg_weight_4_3), .reg_partial_sum(spare_reg_psum_4_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_4( .activation_in(spare_reg_activation_4_3), .weight_in(spare_reg_weight_3_4), .partial_sum_in(spare_reg_psum_3_4), .reg_activation(spare_reg_activation_4_4), .reg_weight(spare_reg_weight_4_4), .reg_partial_sum(spare_reg_psum_4_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_5( .activation_in(spare_reg_activation_4_4), .weight_in(spare_reg_weight_3_5), .partial_sum_in(spare_reg_psum_3_5), .reg_activation(spare_reg_activation_4_5), .reg_weight(spare_reg_weight_4_5), .reg_partial_sum(spare_reg_psum_4_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_6( .activation_in(spare_reg_activation_4_5), .weight_in(spare_reg_weight_3_6), .partial_sum_in(spare_reg_psum_3_6), .reg_activation(spare_reg_activation_4_6), .reg_weight(spare_reg_weight_4_6), .reg_partial_sum(spare_reg_psum_4_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_7( .activation_in(spare_reg_activation_4_6), .weight_in(spare_reg_weight_3_7), .partial_sum_in(spare_reg_psum_3_7), .reg_activation(spare_reg_activation_4_7), .reg_weight(spare_reg_weight_4_7), .reg_partial_sum(spare_reg_psum_4_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_8( .activation_in(spare_reg_activation_4_7), .weight_in(spare_reg_weight_3_8), .partial_sum_in(spare_reg_psum_3_8), .reg_activation(spare_reg_activation_4_8), .reg_weight(spare_reg_weight_4_8), .reg_partial_sum(spare_reg_psum_4_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_9( .activation_in(spare_reg_activation_4_8), .weight_in(spare_reg_weight_3_9), .partial_sum_in(spare_reg_psum_3_9), .reg_activation(spare_reg_activation_4_9), .reg_weight(spare_reg_weight_4_9), .reg_partial_sum(spare_reg_psum_4_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_10( .activation_in(spare_reg_activation_4_9), .weight_in(spare_reg_weight_3_10), .partial_sum_in(spare_reg_psum_3_10), .reg_activation(spare_reg_activation_4_10), .reg_weight(spare_reg_weight_4_10), .reg_partial_sum(spare_reg_psum_4_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_11( .activation_in(spare_reg_activation_4_10), .weight_in(spare_reg_weight_3_11), .partial_sum_in(spare_reg_psum_3_11), .reg_activation(spare_reg_activation_4_11), .reg_weight(spare_reg_weight_4_11), .reg_partial_sum(spare_reg_psum_4_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_12( .activation_in(spare_reg_activation_4_11), .weight_in(spare_reg_weight_3_12), .partial_sum_in(spare_reg_psum_3_12), .reg_activation(spare_reg_activation_4_12), .reg_weight(spare_reg_weight_4_12), .reg_partial_sum(spare_reg_psum_4_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_13( .activation_in(spare_reg_activation_4_12), .weight_in(spare_reg_weight_3_13), .partial_sum_in(spare_reg_psum_3_13), .reg_activation(spare_reg_activation_4_13), .reg_weight(spare_reg_weight_4_13), .reg_partial_sum(spare_reg_psum_4_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_14( .activation_in(spare_reg_activation_4_13), .weight_in(spare_reg_weight_3_14), .partial_sum_in(spare_reg_psum_3_14), .reg_activation(spare_reg_activation_4_14), .reg_weight(spare_reg_weight_4_14), .reg_partial_sum(spare_reg_psum_4_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_15( .activation_in(spare_reg_activation_4_14), .weight_in(spare_reg_weight_3_15), .partial_sum_in(spare_reg_psum_3_15), .reg_activation(spare_reg_activation_4_15), .reg_weight(spare_reg_weight_4_15), .reg_partial_sum(spare_reg_psum_4_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_16( .activation_in(spare_reg_activation_4_15), .weight_in(spare_reg_weight_3_16), .partial_sum_in(spare_reg_psum_3_16), .reg_activation(spare_reg_activation_4_16), .reg_weight(spare_reg_weight_4_16), .reg_partial_sum(spare_reg_psum_4_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_17( .activation_in(spare_reg_activation_4_16), .weight_in(spare_reg_weight_3_17), .partial_sum_in(spare_reg_psum_3_17), .reg_activation(spare_reg_activation_4_17), .reg_weight(spare_reg_weight_4_17), .reg_partial_sum(spare_reg_psum_4_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_18( .activation_in(spare_reg_activation_4_17), .weight_in(spare_reg_weight_3_18), .partial_sum_in(spare_reg_psum_3_18), .reg_activation(spare_reg_activation_4_18), .reg_weight(spare_reg_weight_4_18), .reg_partial_sum(spare_reg_psum_4_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_19( .activation_in(spare_reg_activation_4_18), .weight_in(spare_reg_weight_3_19), .partial_sum_in(spare_reg_psum_3_19), .reg_activation(spare_reg_activation_4_19), .reg_weight(spare_reg_weight_4_19), .reg_partial_sum(spare_reg_psum_4_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_20( .activation_in(spare_reg_activation_4_19), .weight_in(spare_reg_weight_3_20), .partial_sum_in(spare_reg_psum_3_20), .reg_activation(spare_reg_activation_4_20), .reg_weight(spare_reg_weight_4_20), .reg_partial_sum(spare_reg_psum_4_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_21( .activation_in(spare_reg_activation_4_20), .weight_in(spare_reg_weight_3_21), .partial_sum_in(spare_reg_psum_3_21), .reg_activation(spare_reg_activation_4_21), .reg_weight(spare_reg_weight_4_21), .reg_partial_sum(spare_reg_psum_4_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_22( .activation_in(spare_reg_activation_4_21), .weight_in(spare_reg_weight_3_22), .partial_sum_in(spare_reg_psum_3_22), .reg_activation(spare_reg_activation_4_22), .reg_weight(spare_reg_weight_4_22), .reg_partial_sum(spare_reg_psum_4_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_23( .activation_in(spare_reg_activation_4_22), .weight_in(spare_reg_weight_3_23), .partial_sum_in(spare_reg_psum_3_23), .reg_activation(spare_reg_activation_4_23), .reg_weight(spare_reg_weight_4_23), .reg_partial_sum(spare_reg_psum_4_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_24( .activation_in(spare_reg_activation_4_23), .weight_in(spare_reg_weight_3_24), .partial_sum_in(spare_reg_psum_3_24), .reg_activation(spare_reg_activation_4_24), .reg_weight(spare_reg_weight_4_24), .reg_partial_sum(spare_reg_psum_4_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_25( .activation_in(spare_reg_activation_4_24), .weight_in(spare_reg_weight_3_25), .partial_sum_in(spare_reg_psum_3_25), .reg_activation(spare_reg_activation_4_25), .reg_weight(spare_reg_weight_4_25), .reg_partial_sum(spare_reg_psum_4_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_26( .activation_in(spare_reg_activation_4_25), .weight_in(spare_reg_weight_3_26), .partial_sum_in(spare_reg_psum_3_26), .reg_activation(spare_reg_activation_4_26), .reg_weight(spare_reg_weight_4_26), .reg_partial_sum(spare_reg_psum_4_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_27( .activation_in(spare_reg_activation_4_26), .weight_in(spare_reg_weight_3_27), .partial_sum_in(spare_reg_psum_3_27), .reg_activation(spare_reg_activation_4_27), .reg_weight(spare_reg_weight_4_27), .reg_partial_sum(spare_reg_psum_4_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_28( .activation_in(spare_reg_activation_4_27), .weight_in(spare_reg_weight_3_28), .partial_sum_in(spare_reg_psum_3_28), .reg_activation(spare_reg_activation_4_28), .reg_weight(spare_reg_weight_4_28), .reg_partial_sum(spare_reg_psum_4_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_29( .activation_in(spare_reg_activation_4_28), .weight_in(spare_reg_weight_3_29), .partial_sum_in(spare_reg_psum_3_29), .reg_activation(spare_reg_activation_4_29), .reg_weight(spare_reg_weight_4_29), .reg_partial_sum(spare_reg_psum_4_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_30( .activation_in(spare_reg_activation_4_29), .weight_in(spare_reg_weight_3_30), .partial_sum_in(spare_reg_psum_3_30), .reg_activation(spare_reg_activation_4_30), .reg_weight(spare_reg_weight_4_30), .reg_partial_sum(spare_reg_psum_4_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X4_31( .activation_in(spare_reg_activation_4_30), .weight_in(spare_reg_weight_3_31), .partial_sum_in(spare_reg_psum_3_31), .reg_weight(spare_reg_weight_4_31), .reg_partial_sum(spare_reg_psum_4_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_0( .activation_in(in_activation_5), .weight_in(spare_reg_weight_4_0), .partial_sum_in(spare_reg_psum_4_0), .reg_activation(spare_reg_activation_5_0), .reg_weight(spare_reg_weight_5_0), .reg_partial_sum(spare_reg_psum_5_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_1( .activation_in(spare_reg_activation_5_0), .weight_in(spare_reg_weight_4_1), .partial_sum_in(spare_reg_psum_4_1), .reg_activation(spare_reg_activation_5_1), .reg_weight(spare_reg_weight_5_1), .reg_partial_sum(spare_reg_psum_5_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_2( .activation_in(spare_reg_activation_5_1), .weight_in(spare_reg_weight_4_2), .partial_sum_in(spare_reg_psum_4_2), .reg_activation(spare_reg_activation_5_2), .reg_weight(spare_reg_weight_5_2), .reg_partial_sum(spare_reg_psum_5_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_3( .activation_in(spare_reg_activation_5_2), .weight_in(spare_reg_weight_4_3), .partial_sum_in(spare_reg_psum_4_3), .reg_activation(spare_reg_activation_5_3), .reg_weight(spare_reg_weight_5_3), .reg_partial_sum(spare_reg_psum_5_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_4( .activation_in(spare_reg_activation_5_3), .weight_in(spare_reg_weight_4_4), .partial_sum_in(spare_reg_psum_4_4), .reg_activation(spare_reg_activation_5_4), .reg_weight(spare_reg_weight_5_4), .reg_partial_sum(spare_reg_psum_5_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_5( .activation_in(spare_reg_activation_5_4), .weight_in(spare_reg_weight_4_5), .partial_sum_in(spare_reg_psum_4_5), .reg_activation(spare_reg_activation_5_5), .reg_weight(spare_reg_weight_5_5), .reg_partial_sum(spare_reg_psum_5_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_6( .activation_in(spare_reg_activation_5_5), .weight_in(spare_reg_weight_4_6), .partial_sum_in(spare_reg_psum_4_6), .reg_activation(spare_reg_activation_5_6), .reg_weight(spare_reg_weight_5_6), .reg_partial_sum(spare_reg_psum_5_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_7( .activation_in(spare_reg_activation_5_6), .weight_in(spare_reg_weight_4_7), .partial_sum_in(spare_reg_psum_4_7), .reg_activation(spare_reg_activation_5_7), .reg_weight(spare_reg_weight_5_7), .reg_partial_sum(spare_reg_psum_5_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_8( .activation_in(spare_reg_activation_5_7), .weight_in(spare_reg_weight_4_8), .partial_sum_in(spare_reg_psum_4_8), .reg_activation(spare_reg_activation_5_8), .reg_weight(spare_reg_weight_5_8), .reg_partial_sum(spare_reg_psum_5_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_9( .activation_in(spare_reg_activation_5_8), .weight_in(spare_reg_weight_4_9), .partial_sum_in(spare_reg_psum_4_9), .reg_activation(spare_reg_activation_5_9), .reg_weight(spare_reg_weight_5_9), .reg_partial_sum(spare_reg_psum_5_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_10( .activation_in(spare_reg_activation_5_9), .weight_in(spare_reg_weight_4_10), .partial_sum_in(spare_reg_psum_4_10), .reg_activation(spare_reg_activation_5_10), .reg_weight(spare_reg_weight_5_10), .reg_partial_sum(spare_reg_psum_5_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_11( .activation_in(spare_reg_activation_5_10), .weight_in(spare_reg_weight_4_11), .partial_sum_in(spare_reg_psum_4_11), .reg_activation(spare_reg_activation_5_11), .reg_weight(spare_reg_weight_5_11), .reg_partial_sum(spare_reg_psum_5_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_12( .activation_in(spare_reg_activation_5_11), .weight_in(spare_reg_weight_4_12), .partial_sum_in(spare_reg_psum_4_12), .reg_activation(spare_reg_activation_5_12), .reg_weight(spare_reg_weight_5_12), .reg_partial_sum(spare_reg_psum_5_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_13( .activation_in(spare_reg_activation_5_12), .weight_in(spare_reg_weight_4_13), .partial_sum_in(spare_reg_psum_4_13), .reg_activation(spare_reg_activation_5_13), .reg_weight(spare_reg_weight_5_13), .reg_partial_sum(spare_reg_psum_5_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_14( .activation_in(spare_reg_activation_5_13), .weight_in(spare_reg_weight_4_14), .partial_sum_in(spare_reg_psum_4_14), .reg_activation(spare_reg_activation_5_14), .reg_weight(spare_reg_weight_5_14), .reg_partial_sum(spare_reg_psum_5_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_15( .activation_in(spare_reg_activation_5_14), .weight_in(spare_reg_weight_4_15), .partial_sum_in(spare_reg_psum_4_15), .reg_activation(spare_reg_activation_5_15), .reg_weight(spare_reg_weight_5_15), .reg_partial_sum(spare_reg_psum_5_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_16( .activation_in(spare_reg_activation_5_15), .weight_in(spare_reg_weight_4_16), .partial_sum_in(spare_reg_psum_4_16), .reg_activation(spare_reg_activation_5_16), .reg_weight(spare_reg_weight_5_16), .reg_partial_sum(spare_reg_psum_5_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_17( .activation_in(spare_reg_activation_5_16), .weight_in(spare_reg_weight_4_17), .partial_sum_in(spare_reg_psum_4_17), .reg_activation(spare_reg_activation_5_17), .reg_weight(spare_reg_weight_5_17), .reg_partial_sum(spare_reg_psum_5_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_18( .activation_in(spare_reg_activation_5_17), .weight_in(spare_reg_weight_4_18), .partial_sum_in(spare_reg_psum_4_18), .reg_activation(spare_reg_activation_5_18), .reg_weight(spare_reg_weight_5_18), .reg_partial_sum(spare_reg_psum_5_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_19( .activation_in(spare_reg_activation_5_18), .weight_in(spare_reg_weight_4_19), .partial_sum_in(spare_reg_psum_4_19), .reg_activation(spare_reg_activation_5_19), .reg_weight(spare_reg_weight_5_19), .reg_partial_sum(spare_reg_psum_5_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_20( .activation_in(spare_reg_activation_5_19), .weight_in(spare_reg_weight_4_20), .partial_sum_in(spare_reg_psum_4_20), .reg_activation(spare_reg_activation_5_20), .reg_weight(spare_reg_weight_5_20), .reg_partial_sum(spare_reg_psum_5_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_21( .activation_in(spare_reg_activation_5_20), .weight_in(spare_reg_weight_4_21), .partial_sum_in(spare_reg_psum_4_21), .reg_activation(spare_reg_activation_5_21), .reg_weight(spare_reg_weight_5_21), .reg_partial_sum(spare_reg_psum_5_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_22( .activation_in(spare_reg_activation_5_21), .weight_in(spare_reg_weight_4_22), .partial_sum_in(spare_reg_psum_4_22), .reg_activation(spare_reg_activation_5_22), .reg_weight(spare_reg_weight_5_22), .reg_partial_sum(spare_reg_psum_5_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_23( .activation_in(spare_reg_activation_5_22), .weight_in(spare_reg_weight_4_23), .partial_sum_in(spare_reg_psum_4_23), .reg_activation(spare_reg_activation_5_23), .reg_weight(spare_reg_weight_5_23), .reg_partial_sum(spare_reg_psum_5_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_24( .activation_in(spare_reg_activation_5_23), .weight_in(spare_reg_weight_4_24), .partial_sum_in(spare_reg_psum_4_24), .reg_activation(spare_reg_activation_5_24), .reg_weight(spare_reg_weight_5_24), .reg_partial_sum(spare_reg_psum_5_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_25( .activation_in(spare_reg_activation_5_24), .weight_in(spare_reg_weight_4_25), .partial_sum_in(spare_reg_psum_4_25), .reg_activation(spare_reg_activation_5_25), .reg_weight(spare_reg_weight_5_25), .reg_partial_sum(spare_reg_psum_5_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_26( .activation_in(spare_reg_activation_5_25), .weight_in(spare_reg_weight_4_26), .partial_sum_in(spare_reg_psum_4_26), .reg_activation(spare_reg_activation_5_26), .reg_weight(spare_reg_weight_5_26), .reg_partial_sum(spare_reg_psum_5_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_27( .activation_in(spare_reg_activation_5_26), .weight_in(spare_reg_weight_4_27), .partial_sum_in(spare_reg_psum_4_27), .reg_activation(spare_reg_activation_5_27), .reg_weight(spare_reg_weight_5_27), .reg_partial_sum(spare_reg_psum_5_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_28( .activation_in(spare_reg_activation_5_27), .weight_in(spare_reg_weight_4_28), .partial_sum_in(spare_reg_psum_4_28), .reg_activation(spare_reg_activation_5_28), .reg_weight(spare_reg_weight_5_28), .reg_partial_sum(spare_reg_psum_5_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_29( .activation_in(spare_reg_activation_5_28), .weight_in(spare_reg_weight_4_29), .partial_sum_in(spare_reg_psum_4_29), .reg_activation(spare_reg_activation_5_29), .reg_weight(spare_reg_weight_5_29), .reg_partial_sum(spare_reg_psum_5_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_30( .activation_in(spare_reg_activation_5_29), .weight_in(spare_reg_weight_4_30), .partial_sum_in(spare_reg_psum_4_30), .reg_activation(spare_reg_activation_5_30), .reg_weight(spare_reg_weight_5_30), .reg_partial_sum(spare_reg_psum_5_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X5_31( .activation_in(spare_reg_activation_5_30), .weight_in(spare_reg_weight_4_31), .partial_sum_in(spare_reg_psum_4_31), .reg_weight(spare_reg_weight_5_31), .reg_partial_sum(spare_reg_psum_5_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_0( .activation_in(in_activation_6), .weight_in(spare_reg_weight_5_0), .partial_sum_in(spare_reg_psum_5_0), .reg_activation(spare_reg_activation_6_0), .reg_weight(spare_reg_weight_6_0), .reg_partial_sum(spare_reg_psum_6_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_1( .activation_in(spare_reg_activation_6_0), .weight_in(spare_reg_weight_5_1), .partial_sum_in(spare_reg_psum_5_1), .reg_activation(spare_reg_activation_6_1), .reg_weight(spare_reg_weight_6_1), .reg_partial_sum(spare_reg_psum_6_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_2( .activation_in(spare_reg_activation_6_1), .weight_in(spare_reg_weight_5_2), .partial_sum_in(spare_reg_psum_5_2), .reg_activation(spare_reg_activation_6_2), .reg_weight(spare_reg_weight_6_2), .reg_partial_sum(spare_reg_psum_6_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_3( .activation_in(spare_reg_activation_6_2), .weight_in(spare_reg_weight_5_3), .partial_sum_in(spare_reg_psum_5_3), .reg_activation(spare_reg_activation_6_3), .reg_weight(spare_reg_weight_6_3), .reg_partial_sum(spare_reg_psum_6_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_4( .activation_in(spare_reg_activation_6_3), .weight_in(spare_reg_weight_5_4), .partial_sum_in(spare_reg_psum_5_4), .reg_activation(spare_reg_activation_6_4), .reg_weight(spare_reg_weight_6_4), .reg_partial_sum(spare_reg_psum_6_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_5( .activation_in(spare_reg_activation_6_4), .weight_in(spare_reg_weight_5_5), .partial_sum_in(spare_reg_psum_5_5), .reg_activation(spare_reg_activation_6_5), .reg_weight(spare_reg_weight_6_5), .reg_partial_sum(spare_reg_psum_6_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_6( .activation_in(spare_reg_activation_6_5), .weight_in(spare_reg_weight_5_6), .partial_sum_in(spare_reg_psum_5_6), .reg_activation(spare_reg_activation_6_6), .reg_weight(spare_reg_weight_6_6), .reg_partial_sum(spare_reg_psum_6_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_7( .activation_in(spare_reg_activation_6_6), .weight_in(spare_reg_weight_5_7), .partial_sum_in(spare_reg_psum_5_7), .reg_activation(spare_reg_activation_6_7), .reg_weight(spare_reg_weight_6_7), .reg_partial_sum(spare_reg_psum_6_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_8( .activation_in(spare_reg_activation_6_7), .weight_in(spare_reg_weight_5_8), .partial_sum_in(spare_reg_psum_5_8), .reg_activation(spare_reg_activation_6_8), .reg_weight(spare_reg_weight_6_8), .reg_partial_sum(spare_reg_psum_6_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_9( .activation_in(spare_reg_activation_6_8), .weight_in(spare_reg_weight_5_9), .partial_sum_in(spare_reg_psum_5_9), .reg_activation(spare_reg_activation_6_9), .reg_weight(spare_reg_weight_6_9), .reg_partial_sum(spare_reg_psum_6_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_10( .activation_in(spare_reg_activation_6_9), .weight_in(spare_reg_weight_5_10), .partial_sum_in(spare_reg_psum_5_10), .reg_activation(spare_reg_activation_6_10), .reg_weight(spare_reg_weight_6_10), .reg_partial_sum(spare_reg_psum_6_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_11( .activation_in(spare_reg_activation_6_10), .weight_in(spare_reg_weight_5_11), .partial_sum_in(spare_reg_psum_5_11), .reg_activation(spare_reg_activation_6_11), .reg_weight(spare_reg_weight_6_11), .reg_partial_sum(spare_reg_psum_6_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_12( .activation_in(spare_reg_activation_6_11), .weight_in(spare_reg_weight_5_12), .partial_sum_in(spare_reg_psum_5_12), .reg_activation(spare_reg_activation_6_12), .reg_weight(spare_reg_weight_6_12), .reg_partial_sum(spare_reg_psum_6_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_13( .activation_in(spare_reg_activation_6_12), .weight_in(spare_reg_weight_5_13), .partial_sum_in(spare_reg_psum_5_13), .reg_activation(spare_reg_activation_6_13), .reg_weight(spare_reg_weight_6_13), .reg_partial_sum(spare_reg_psum_6_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_14( .activation_in(spare_reg_activation_6_13), .weight_in(spare_reg_weight_5_14), .partial_sum_in(spare_reg_psum_5_14), .reg_activation(spare_reg_activation_6_14), .reg_weight(spare_reg_weight_6_14), .reg_partial_sum(spare_reg_psum_6_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_15( .activation_in(spare_reg_activation_6_14), .weight_in(spare_reg_weight_5_15), .partial_sum_in(spare_reg_psum_5_15), .reg_activation(spare_reg_activation_6_15), .reg_weight(spare_reg_weight_6_15), .reg_partial_sum(spare_reg_psum_6_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_16( .activation_in(spare_reg_activation_6_15), .weight_in(spare_reg_weight_5_16), .partial_sum_in(spare_reg_psum_5_16), .reg_activation(spare_reg_activation_6_16), .reg_weight(spare_reg_weight_6_16), .reg_partial_sum(spare_reg_psum_6_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_17( .activation_in(spare_reg_activation_6_16), .weight_in(spare_reg_weight_5_17), .partial_sum_in(spare_reg_psum_5_17), .reg_activation(spare_reg_activation_6_17), .reg_weight(spare_reg_weight_6_17), .reg_partial_sum(spare_reg_psum_6_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_18( .activation_in(spare_reg_activation_6_17), .weight_in(spare_reg_weight_5_18), .partial_sum_in(spare_reg_psum_5_18), .reg_activation(spare_reg_activation_6_18), .reg_weight(spare_reg_weight_6_18), .reg_partial_sum(spare_reg_psum_6_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_19( .activation_in(spare_reg_activation_6_18), .weight_in(spare_reg_weight_5_19), .partial_sum_in(spare_reg_psum_5_19), .reg_activation(spare_reg_activation_6_19), .reg_weight(spare_reg_weight_6_19), .reg_partial_sum(spare_reg_psum_6_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_20( .activation_in(spare_reg_activation_6_19), .weight_in(spare_reg_weight_5_20), .partial_sum_in(spare_reg_psum_5_20), .reg_activation(spare_reg_activation_6_20), .reg_weight(spare_reg_weight_6_20), .reg_partial_sum(spare_reg_psum_6_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_21( .activation_in(spare_reg_activation_6_20), .weight_in(spare_reg_weight_5_21), .partial_sum_in(spare_reg_psum_5_21), .reg_activation(spare_reg_activation_6_21), .reg_weight(spare_reg_weight_6_21), .reg_partial_sum(spare_reg_psum_6_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_22( .activation_in(spare_reg_activation_6_21), .weight_in(spare_reg_weight_5_22), .partial_sum_in(spare_reg_psum_5_22), .reg_activation(spare_reg_activation_6_22), .reg_weight(spare_reg_weight_6_22), .reg_partial_sum(spare_reg_psum_6_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_23( .activation_in(spare_reg_activation_6_22), .weight_in(spare_reg_weight_5_23), .partial_sum_in(spare_reg_psum_5_23), .reg_activation(spare_reg_activation_6_23), .reg_weight(spare_reg_weight_6_23), .reg_partial_sum(spare_reg_psum_6_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_24( .activation_in(spare_reg_activation_6_23), .weight_in(spare_reg_weight_5_24), .partial_sum_in(spare_reg_psum_5_24), .reg_activation(spare_reg_activation_6_24), .reg_weight(spare_reg_weight_6_24), .reg_partial_sum(spare_reg_psum_6_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_25( .activation_in(spare_reg_activation_6_24), .weight_in(spare_reg_weight_5_25), .partial_sum_in(spare_reg_psum_5_25), .reg_activation(spare_reg_activation_6_25), .reg_weight(spare_reg_weight_6_25), .reg_partial_sum(spare_reg_psum_6_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_26( .activation_in(spare_reg_activation_6_25), .weight_in(spare_reg_weight_5_26), .partial_sum_in(spare_reg_psum_5_26), .reg_activation(spare_reg_activation_6_26), .reg_weight(spare_reg_weight_6_26), .reg_partial_sum(spare_reg_psum_6_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_27( .activation_in(spare_reg_activation_6_26), .weight_in(spare_reg_weight_5_27), .partial_sum_in(spare_reg_psum_5_27), .reg_activation(spare_reg_activation_6_27), .reg_weight(spare_reg_weight_6_27), .reg_partial_sum(spare_reg_psum_6_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_28( .activation_in(spare_reg_activation_6_27), .weight_in(spare_reg_weight_5_28), .partial_sum_in(spare_reg_psum_5_28), .reg_activation(spare_reg_activation_6_28), .reg_weight(spare_reg_weight_6_28), .reg_partial_sum(spare_reg_psum_6_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_29( .activation_in(spare_reg_activation_6_28), .weight_in(spare_reg_weight_5_29), .partial_sum_in(spare_reg_psum_5_29), .reg_activation(spare_reg_activation_6_29), .reg_weight(spare_reg_weight_6_29), .reg_partial_sum(spare_reg_psum_6_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_30( .activation_in(spare_reg_activation_6_29), .weight_in(spare_reg_weight_5_30), .partial_sum_in(spare_reg_psum_5_30), .reg_activation(spare_reg_activation_6_30), .reg_weight(spare_reg_weight_6_30), .reg_partial_sum(spare_reg_psum_6_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X6_31( .activation_in(spare_reg_activation_6_30), .weight_in(spare_reg_weight_5_31), .partial_sum_in(spare_reg_psum_5_31), .reg_weight(spare_reg_weight_6_31), .reg_partial_sum(spare_reg_psum_6_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_0( .activation_in(in_activation_7), .weight_in(spare_reg_weight_6_0), .partial_sum_in(spare_reg_psum_6_0), .reg_activation(spare_reg_activation_7_0), .reg_weight(spare_reg_weight_7_0), .reg_partial_sum(spare_reg_psum_7_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_1( .activation_in(spare_reg_activation_7_0), .weight_in(spare_reg_weight_6_1), .partial_sum_in(spare_reg_psum_6_1), .reg_activation(spare_reg_activation_7_1), .reg_weight(spare_reg_weight_7_1), .reg_partial_sum(spare_reg_psum_7_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_2( .activation_in(spare_reg_activation_7_1), .weight_in(spare_reg_weight_6_2), .partial_sum_in(spare_reg_psum_6_2), .reg_activation(spare_reg_activation_7_2), .reg_weight(spare_reg_weight_7_2), .reg_partial_sum(spare_reg_psum_7_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_3( .activation_in(spare_reg_activation_7_2), .weight_in(spare_reg_weight_6_3), .partial_sum_in(spare_reg_psum_6_3), .reg_activation(spare_reg_activation_7_3), .reg_weight(spare_reg_weight_7_3), .reg_partial_sum(spare_reg_psum_7_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_4( .activation_in(spare_reg_activation_7_3), .weight_in(spare_reg_weight_6_4), .partial_sum_in(spare_reg_psum_6_4), .reg_activation(spare_reg_activation_7_4), .reg_weight(spare_reg_weight_7_4), .reg_partial_sum(spare_reg_psum_7_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_5( .activation_in(spare_reg_activation_7_4), .weight_in(spare_reg_weight_6_5), .partial_sum_in(spare_reg_psum_6_5), .reg_activation(spare_reg_activation_7_5), .reg_weight(spare_reg_weight_7_5), .reg_partial_sum(spare_reg_psum_7_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_6( .activation_in(spare_reg_activation_7_5), .weight_in(spare_reg_weight_6_6), .partial_sum_in(spare_reg_psum_6_6), .reg_activation(spare_reg_activation_7_6), .reg_weight(spare_reg_weight_7_6), .reg_partial_sum(spare_reg_psum_7_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_7( .activation_in(spare_reg_activation_7_6), .weight_in(spare_reg_weight_6_7), .partial_sum_in(spare_reg_psum_6_7), .reg_activation(spare_reg_activation_7_7), .reg_weight(spare_reg_weight_7_7), .reg_partial_sum(spare_reg_psum_7_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_8( .activation_in(spare_reg_activation_7_7), .weight_in(spare_reg_weight_6_8), .partial_sum_in(spare_reg_psum_6_8), .reg_activation(spare_reg_activation_7_8), .reg_weight(spare_reg_weight_7_8), .reg_partial_sum(spare_reg_psum_7_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_9( .activation_in(spare_reg_activation_7_8), .weight_in(spare_reg_weight_6_9), .partial_sum_in(spare_reg_psum_6_9), .reg_activation(spare_reg_activation_7_9), .reg_weight(spare_reg_weight_7_9), .reg_partial_sum(spare_reg_psum_7_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_10( .activation_in(spare_reg_activation_7_9), .weight_in(spare_reg_weight_6_10), .partial_sum_in(spare_reg_psum_6_10), .reg_activation(spare_reg_activation_7_10), .reg_weight(spare_reg_weight_7_10), .reg_partial_sum(spare_reg_psum_7_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_11( .activation_in(spare_reg_activation_7_10), .weight_in(spare_reg_weight_6_11), .partial_sum_in(spare_reg_psum_6_11), .reg_activation(spare_reg_activation_7_11), .reg_weight(spare_reg_weight_7_11), .reg_partial_sum(spare_reg_psum_7_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_12( .activation_in(spare_reg_activation_7_11), .weight_in(spare_reg_weight_6_12), .partial_sum_in(spare_reg_psum_6_12), .reg_activation(spare_reg_activation_7_12), .reg_weight(spare_reg_weight_7_12), .reg_partial_sum(spare_reg_psum_7_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_13( .activation_in(spare_reg_activation_7_12), .weight_in(spare_reg_weight_6_13), .partial_sum_in(spare_reg_psum_6_13), .reg_activation(spare_reg_activation_7_13), .reg_weight(spare_reg_weight_7_13), .reg_partial_sum(spare_reg_psum_7_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_14( .activation_in(spare_reg_activation_7_13), .weight_in(spare_reg_weight_6_14), .partial_sum_in(spare_reg_psum_6_14), .reg_activation(spare_reg_activation_7_14), .reg_weight(spare_reg_weight_7_14), .reg_partial_sum(spare_reg_psum_7_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_15( .activation_in(spare_reg_activation_7_14), .weight_in(spare_reg_weight_6_15), .partial_sum_in(spare_reg_psum_6_15), .reg_activation(spare_reg_activation_7_15), .reg_weight(spare_reg_weight_7_15), .reg_partial_sum(spare_reg_psum_7_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_16( .activation_in(spare_reg_activation_7_15), .weight_in(spare_reg_weight_6_16), .partial_sum_in(spare_reg_psum_6_16), .reg_activation(spare_reg_activation_7_16), .reg_weight(spare_reg_weight_7_16), .reg_partial_sum(spare_reg_psum_7_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_17( .activation_in(spare_reg_activation_7_16), .weight_in(spare_reg_weight_6_17), .partial_sum_in(spare_reg_psum_6_17), .reg_activation(spare_reg_activation_7_17), .reg_weight(spare_reg_weight_7_17), .reg_partial_sum(spare_reg_psum_7_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_18( .activation_in(spare_reg_activation_7_17), .weight_in(spare_reg_weight_6_18), .partial_sum_in(spare_reg_psum_6_18), .reg_activation(spare_reg_activation_7_18), .reg_weight(spare_reg_weight_7_18), .reg_partial_sum(spare_reg_psum_7_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_19( .activation_in(spare_reg_activation_7_18), .weight_in(spare_reg_weight_6_19), .partial_sum_in(spare_reg_psum_6_19), .reg_activation(spare_reg_activation_7_19), .reg_weight(spare_reg_weight_7_19), .reg_partial_sum(spare_reg_psum_7_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_20( .activation_in(spare_reg_activation_7_19), .weight_in(spare_reg_weight_6_20), .partial_sum_in(spare_reg_psum_6_20), .reg_activation(spare_reg_activation_7_20), .reg_weight(spare_reg_weight_7_20), .reg_partial_sum(spare_reg_psum_7_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_21( .activation_in(spare_reg_activation_7_20), .weight_in(spare_reg_weight_6_21), .partial_sum_in(spare_reg_psum_6_21), .reg_activation(spare_reg_activation_7_21), .reg_weight(spare_reg_weight_7_21), .reg_partial_sum(spare_reg_psum_7_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_22( .activation_in(spare_reg_activation_7_21), .weight_in(spare_reg_weight_6_22), .partial_sum_in(spare_reg_psum_6_22), .reg_activation(spare_reg_activation_7_22), .reg_weight(spare_reg_weight_7_22), .reg_partial_sum(spare_reg_psum_7_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_23( .activation_in(spare_reg_activation_7_22), .weight_in(spare_reg_weight_6_23), .partial_sum_in(spare_reg_psum_6_23), .reg_activation(spare_reg_activation_7_23), .reg_weight(spare_reg_weight_7_23), .reg_partial_sum(spare_reg_psum_7_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_24( .activation_in(spare_reg_activation_7_23), .weight_in(spare_reg_weight_6_24), .partial_sum_in(spare_reg_psum_6_24), .reg_activation(spare_reg_activation_7_24), .reg_weight(spare_reg_weight_7_24), .reg_partial_sum(spare_reg_psum_7_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_25( .activation_in(spare_reg_activation_7_24), .weight_in(spare_reg_weight_6_25), .partial_sum_in(spare_reg_psum_6_25), .reg_activation(spare_reg_activation_7_25), .reg_weight(spare_reg_weight_7_25), .reg_partial_sum(spare_reg_psum_7_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_26( .activation_in(spare_reg_activation_7_25), .weight_in(spare_reg_weight_6_26), .partial_sum_in(spare_reg_psum_6_26), .reg_activation(spare_reg_activation_7_26), .reg_weight(spare_reg_weight_7_26), .reg_partial_sum(spare_reg_psum_7_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_27( .activation_in(spare_reg_activation_7_26), .weight_in(spare_reg_weight_6_27), .partial_sum_in(spare_reg_psum_6_27), .reg_activation(spare_reg_activation_7_27), .reg_weight(spare_reg_weight_7_27), .reg_partial_sum(spare_reg_psum_7_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_28( .activation_in(spare_reg_activation_7_27), .weight_in(spare_reg_weight_6_28), .partial_sum_in(spare_reg_psum_6_28), .reg_activation(spare_reg_activation_7_28), .reg_weight(spare_reg_weight_7_28), .reg_partial_sum(spare_reg_psum_7_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_29( .activation_in(spare_reg_activation_7_28), .weight_in(spare_reg_weight_6_29), .partial_sum_in(spare_reg_psum_6_29), .reg_activation(spare_reg_activation_7_29), .reg_weight(spare_reg_weight_7_29), .reg_partial_sum(spare_reg_psum_7_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_30( .activation_in(spare_reg_activation_7_29), .weight_in(spare_reg_weight_6_30), .partial_sum_in(spare_reg_psum_6_30), .reg_activation(spare_reg_activation_7_30), .reg_weight(spare_reg_weight_7_30), .reg_partial_sum(spare_reg_psum_7_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X7_31( .activation_in(spare_reg_activation_7_30), .weight_in(spare_reg_weight_6_31), .partial_sum_in(spare_reg_psum_6_31), .reg_weight(spare_reg_weight_7_31), .reg_partial_sum(spare_reg_psum_7_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_0( .activation_in(in_activation_8), .weight_in(spare_reg_weight_7_0), .partial_sum_in(spare_reg_psum_7_0), .reg_activation(spare_reg_activation_8_0), .reg_weight(spare_reg_weight_8_0), .reg_partial_sum(spare_reg_psum_8_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_1( .activation_in(spare_reg_activation_8_0), .weight_in(spare_reg_weight_7_1), .partial_sum_in(spare_reg_psum_7_1), .reg_activation(spare_reg_activation_8_1), .reg_weight(spare_reg_weight_8_1), .reg_partial_sum(spare_reg_psum_8_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_2( .activation_in(spare_reg_activation_8_1), .weight_in(spare_reg_weight_7_2), .partial_sum_in(spare_reg_psum_7_2), .reg_activation(spare_reg_activation_8_2), .reg_weight(spare_reg_weight_8_2), .reg_partial_sum(spare_reg_psum_8_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_3( .activation_in(spare_reg_activation_8_2), .weight_in(spare_reg_weight_7_3), .partial_sum_in(spare_reg_psum_7_3), .reg_activation(spare_reg_activation_8_3), .reg_weight(spare_reg_weight_8_3), .reg_partial_sum(spare_reg_psum_8_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_4( .activation_in(spare_reg_activation_8_3), .weight_in(spare_reg_weight_7_4), .partial_sum_in(spare_reg_psum_7_4), .reg_activation(spare_reg_activation_8_4), .reg_weight(spare_reg_weight_8_4), .reg_partial_sum(spare_reg_psum_8_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_5( .activation_in(spare_reg_activation_8_4), .weight_in(spare_reg_weight_7_5), .partial_sum_in(spare_reg_psum_7_5), .reg_activation(spare_reg_activation_8_5), .reg_weight(spare_reg_weight_8_5), .reg_partial_sum(spare_reg_psum_8_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_6( .activation_in(spare_reg_activation_8_5), .weight_in(spare_reg_weight_7_6), .partial_sum_in(spare_reg_psum_7_6), .reg_activation(spare_reg_activation_8_6), .reg_weight(spare_reg_weight_8_6), .reg_partial_sum(spare_reg_psum_8_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_7( .activation_in(spare_reg_activation_8_6), .weight_in(spare_reg_weight_7_7), .partial_sum_in(spare_reg_psum_7_7), .reg_activation(spare_reg_activation_8_7), .reg_weight(spare_reg_weight_8_7), .reg_partial_sum(spare_reg_psum_8_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_8( .activation_in(spare_reg_activation_8_7), .weight_in(spare_reg_weight_7_8), .partial_sum_in(spare_reg_psum_7_8), .reg_activation(spare_reg_activation_8_8), .reg_weight(spare_reg_weight_8_8), .reg_partial_sum(spare_reg_psum_8_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_9( .activation_in(spare_reg_activation_8_8), .weight_in(spare_reg_weight_7_9), .partial_sum_in(spare_reg_psum_7_9), .reg_activation(spare_reg_activation_8_9), .reg_weight(spare_reg_weight_8_9), .reg_partial_sum(spare_reg_psum_8_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_10( .activation_in(spare_reg_activation_8_9), .weight_in(spare_reg_weight_7_10), .partial_sum_in(spare_reg_psum_7_10), .reg_activation(spare_reg_activation_8_10), .reg_weight(spare_reg_weight_8_10), .reg_partial_sum(spare_reg_psum_8_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_11( .activation_in(spare_reg_activation_8_10), .weight_in(spare_reg_weight_7_11), .partial_sum_in(spare_reg_psum_7_11), .reg_activation(spare_reg_activation_8_11), .reg_weight(spare_reg_weight_8_11), .reg_partial_sum(spare_reg_psum_8_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_12( .activation_in(spare_reg_activation_8_11), .weight_in(spare_reg_weight_7_12), .partial_sum_in(spare_reg_psum_7_12), .reg_activation(spare_reg_activation_8_12), .reg_weight(spare_reg_weight_8_12), .reg_partial_sum(spare_reg_psum_8_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_13( .activation_in(spare_reg_activation_8_12), .weight_in(spare_reg_weight_7_13), .partial_sum_in(spare_reg_psum_7_13), .reg_activation(spare_reg_activation_8_13), .reg_weight(spare_reg_weight_8_13), .reg_partial_sum(spare_reg_psum_8_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_14( .activation_in(spare_reg_activation_8_13), .weight_in(spare_reg_weight_7_14), .partial_sum_in(spare_reg_psum_7_14), .reg_activation(spare_reg_activation_8_14), .reg_weight(spare_reg_weight_8_14), .reg_partial_sum(spare_reg_psum_8_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_15( .activation_in(spare_reg_activation_8_14), .weight_in(spare_reg_weight_7_15), .partial_sum_in(spare_reg_psum_7_15), .reg_activation(spare_reg_activation_8_15), .reg_weight(spare_reg_weight_8_15), .reg_partial_sum(spare_reg_psum_8_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_16( .activation_in(spare_reg_activation_8_15), .weight_in(spare_reg_weight_7_16), .partial_sum_in(spare_reg_psum_7_16), .reg_activation(spare_reg_activation_8_16), .reg_weight(spare_reg_weight_8_16), .reg_partial_sum(spare_reg_psum_8_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_17( .activation_in(spare_reg_activation_8_16), .weight_in(spare_reg_weight_7_17), .partial_sum_in(spare_reg_psum_7_17), .reg_activation(spare_reg_activation_8_17), .reg_weight(spare_reg_weight_8_17), .reg_partial_sum(spare_reg_psum_8_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_18( .activation_in(spare_reg_activation_8_17), .weight_in(spare_reg_weight_7_18), .partial_sum_in(spare_reg_psum_7_18), .reg_activation(spare_reg_activation_8_18), .reg_weight(spare_reg_weight_8_18), .reg_partial_sum(spare_reg_psum_8_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_19( .activation_in(spare_reg_activation_8_18), .weight_in(spare_reg_weight_7_19), .partial_sum_in(spare_reg_psum_7_19), .reg_activation(spare_reg_activation_8_19), .reg_weight(spare_reg_weight_8_19), .reg_partial_sum(spare_reg_psum_8_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_20( .activation_in(spare_reg_activation_8_19), .weight_in(spare_reg_weight_7_20), .partial_sum_in(spare_reg_psum_7_20), .reg_activation(spare_reg_activation_8_20), .reg_weight(spare_reg_weight_8_20), .reg_partial_sum(spare_reg_psum_8_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_21( .activation_in(spare_reg_activation_8_20), .weight_in(spare_reg_weight_7_21), .partial_sum_in(spare_reg_psum_7_21), .reg_activation(spare_reg_activation_8_21), .reg_weight(spare_reg_weight_8_21), .reg_partial_sum(spare_reg_psum_8_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_22( .activation_in(spare_reg_activation_8_21), .weight_in(spare_reg_weight_7_22), .partial_sum_in(spare_reg_psum_7_22), .reg_activation(spare_reg_activation_8_22), .reg_weight(spare_reg_weight_8_22), .reg_partial_sum(spare_reg_psum_8_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_23( .activation_in(spare_reg_activation_8_22), .weight_in(spare_reg_weight_7_23), .partial_sum_in(spare_reg_psum_7_23), .reg_activation(spare_reg_activation_8_23), .reg_weight(spare_reg_weight_8_23), .reg_partial_sum(spare_reg_psum_8_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_24( .activation_in(spare_reg_activation_8_23), .weight_in(spare_reg_weight_7_24), .partial_sum_in(spare_reg_psum_7_24), .reg_activation(spare_reg_activation_8_24), .reg_weight(spare_reg_weight_8_24), .reg_partial_sum(spare_reg_psum_8_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_25( .activation_in(spare_reg_activation_8_24), .weight_in(spare_reg_weight_7_25), .partial_sum_in(spare_reg_psum_7_25), .reg_activation(spare_reg_activation_8_25), .reg_weight(spare_reg_weight_8_25), .reg_partial_sum(spare_reg_psum_8_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_26( .activation_in(spare_reg_activation_8_25), .weight_in(spare_reg_weight_7_26), .partial_sum_in(spare_reg_psum_7_26), .reg_activation(spare_reg_activation_8_26), .reg_weight(spare_reg_weight_8_26), .reg_partial_sum(spare_reg_psum_8_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_27( .activation_in(spare_reg_activation_8_26), .weight_in(spare_reg_weight_7_27), .partial_sum_in(spare_reg_psum_7_27), .reg_activation(spare_reg_activation_8_27), .reg_weight(spare_reg_weight_8_27), .reg_partial_sum(spare_reg_psum_8_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_28( .activation_in(spare_reg_activation_8_27), .weight_in(spare_reg_weight_7_28), .partial_sum_in(spare_reg_psum_7_28), .reg_activation(spare_reg_activation_8_28), .reg_weight(spare_reg_weight_8_28), .reg_partial_sum(spare_reg_psum_8_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_29( .activation_in(spare_reg_activation_8_28), .weight_in(spare_reg_weight_7_29), .partial_sum_in(spare_reg_psum_7_29), .reg_activation(spare_reg_activation_8_29), .reg_weight(spare_reg_weight_8_29), .reg_partial_sum(spare_reg_psum_8_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_30( .activation_in(spare_reg_activation_8_29), .weight_in(spare_reg_weight_7_30), .partial_sum_in(spare_reg_psum_7_30), .reg_activation(spare_reg_activation_8_30), .reg_weight(spare_reg_weight_8_30), .reg_partial_sum(spare_reg_psum_8_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X8_31( .activation_in(spare_reg_activation_8_30), .weight_in(spare_reg_weight_7_31), .partial_sum_in(spare_reg_psum_7_31), .reg_weight(spare_reg_weight_8_31), .reg_partial_sum(spare_reg_psum_8_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_0( .activation_in(in_activation_9), .weight_in(spare_reg_weight_8_0), .partial_sum_in(spare_reg_psum_8_0), .reg_activation(spare_reg_activation_9_0), .reg_weight(spare_reg_weight_9_0), .reg_partial_sum(spare_reg_psum_9_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_1( .activation_in(spare_reg_activation_9_0), .weight_in(spare_reg_weight_8_1), .partial_sum_in(spare_reg_psum_8_1), .reg_activation(spare_reg_activation_9_1), .reg_weight(spare_reg_weight_9_1), .reg_partial_sum(spare_reg_psum_9_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_2( .activation_in(spare_reg_activation_9_1), .weight_in(spare_reg_weight_8_2), .partial_sum_in(spare_reg_psum_8_2), .reg_activation(spare_reg_activation_9_2), .reg_weight(spare_reg_weight_9_2), .reg_partial_sum(spare_reg_psum_9_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_3( .activation_in(spare_reg_activation_9_2), .weight_in(spare_reg_weight_8_3), .partial_sum_in(spare_reg_psum_8_3), .reg_activation(spare_reg_activation_9_3), .reg_weight(spare_reg_weight_9_3), .reg_partial_sum(spare_reg_psum_9_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_4( .activation_in(spare_reg_activation_9_3), .weight_in(spare_reg_weight_8_4), .partial_sum_in(spare_reg_psum_8_4), .reg_activation(spare_reg_activation_9_4), .reg_weight(spare_reg_weight_9_4), .reg_partial_sum(spare_reg_psum_9_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_5( .activation_in(spare_reg_activation_9_4), .weight_in(spare_reg_weight_8_5), .partial_sum_in(spare_reg_psum_8_5), .reg_activation(spare_reg_activation_9_5), .reg_weight(spare_reg_weight_9_5), .reg_partial_sum(spare_reg_psum_9_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_6( .activation_in(spare_reg_activation_9_5), .weight_in(spare_reg_weight_8_6), .partial_sum_in(spare_reg_psum_8_6), .reg_activation(spare_reg_activation_9_6), .reg_weight(spare_reg_weight_9_6), .reg_partial_sum(spare_reg_psum_9_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_7( .activation_in(spare_reg_activation_9_6), .weight_in(spare_reg_weight_8_7), .partial_sum_in(spare_reg_psum_8_7), .reg_activation(spare_reg_activation_9_7), .reg_weight(spare_reg_weight_9_7), .reg_partial_sum(spare_reg_psum_9_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_8( .activation_in(spare_reg_activation_9_7), .weight_in(spare_reg_weight_8_8), .partial_sum_in(spare_reg_psum_8_8), .reg_activation(spare_reg_activation_9_8), .reg_weight(spare_reg_weight_9_8), .reg_partial_sum(spare_reg_psum_9_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_9( .activation_in(spare_reg_activation_9_8), .weight_in(spare_reg_weight_8_9), .partial_sum_in(spare_reg_psum_8_9), .reg_activation(spare_reg_activation_9_9), .reg_weight(spare_reg_weight_9_9), .reg_partial_sum(spare_reg_psum_9_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_10( .activation_in(spare_reg_activation_9_9), .weight_in(spare_reg_weight_8_10), .partial_sum_in(spare_reg_psum_8_10), .reg_activation(spare_reg_activation_9_10), .reg_weight(spare_reg_weight_9_10), .reg_partial_sum(spare_reg_psum_9_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_11( .activation_in(spare_reg_activation_9_10), .weight_in(spare_reg_weight_8_11), .partial_sum_in(spare_reg_psum_8_11), .reg_activation(spare_reg_activation_9_11), .reg_weight(spare_reg_weight_9_11), .reg_partial_sum(spare_reg_psum_9_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_12( .activation_in(spare_reg_activation_9_11), .weight_in(spare_reg_weight_8_12), .partial_sum_in(spare_reg_psum_8_12), .reg_activation(spare_reg_activation_9_12), .reg_weight(spare_reg_weight_9_12), .reg_partial_sum(spare_reg_psum_9_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_13( .activation_in(spare_reg_activation_9_12), .weight_in(spare_reg_weight_8_13), .partial_sum_in(spare_reg_psum_8_13), .reg_activation(spare_reg_activation_9_13), .reg_weight(spare_reg_weight_9_13), .reg_partial_sum(spare_reg_psum_9_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_14( .activation_in(spare_reg_activation_9_13), .weight_in(spare_reg_weight_8_14), .partial_sum_in(spare_reg_psum_8_14), .reg_activation(spare_reg_activation_9_14), .reg_weight(spare_reg_weight_9_14), .reg_partial_sum(spare_reg_psum_9_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_15( .activation_in(spare_reg_activation_9_14), .weight_in(spare_reg_weight_8_15), .partial_sum_in(spare_reg_psum_8_15), .reg_activation(spare_reg_activation_9_15), .reg_weight(spare_reg_weight_9_15), .reg_partial_sum(spare_reg_psum_9_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_16( .activation_in(spare_reg_activation_9_15), .weight_in(spare_reg_weight_8_16), .partial_sum_in(spare_reg_psum_8_16), .reg_activation(spare_reg_activation_9_16), .reg_weight(spare_reg_weight_9_16), .reg_partial_sum(spare_reg_psum_9_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_17( .activation_in(spare_reg_activation_9_16), .weight_in(spare_reg_weight_8_17), .partial_sum_in(spare_reg_psum_8_17), .reg_activation(spare_reg_activation_9_17), .reg_weight(spare_reg_weight_9_17), .reg_partial_sum(spare_reg_psum_9_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_18( .activation_in(spare_reg_activation_9_17), .weight_in(spare_reg_weight_8_18), .partial_sum_in(spare_reg_psum_8_18), .reg_activation(spare_reg_activation_9_18), .reg_weight(spare_reg_weight_9_18), .reg_partial_sum(spare_reg_psum_9_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_19( .activation_in(spare_reg_activation_9_18), .weight_in(spare_reg_weight_8_19), .partial_sum_in(spare_reg_psum_8_19), .reg_activation(spare_reg_activation_9_19), .reg_weight(spare_reg_weight_9_19), .reg_partial_sum(spare_reg_psum_9_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_20( .activation_in(spare_reg_activation_9_19), .weight_in(spare_reg_weight_8_20), .partial_sum_in(spare_reg_psum_8_20), .reg_activation(spare_reg_activation_9_20), .reg_weight(spare_reg_weight_9_20), .reg_partial_sum(spare_reg_psum_9_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_21( .activation_in(spare_reg_activation_9_20), .weight_in(spare_reg_weight_8_21), .partial_sum_in(spare_reg_psum_8_21), .reg_activation(spare_reg_activation_9_21), .reg_weight(spare_reg_weight_9_21), .reg_partial_sum(spare_reg_psum_9_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_22( .activation_in(spare_reg_activation_9_21), .weight_in(spare_reg_weight_8_22), .partial_sum_in(spare_reg_psum_8_22), .reg_activation(spare_reg_activation_9_22), .reg_weight(spare_reg_weight_9_22), .reg_partial_sum(spare_reg_psum_9_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_23( .activation_in(spare_reg_activation_9_22), .weight_in(spare_reg_weight_8_23), .partial_sum_in(spare_reg_psum_8_23), .reg_activation(spare_reg_activation_9_23), .reg_weight(spare_reg_weight_9_23), .reg_partial_sum(spare_reg_psum_9_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_24( .activation_in(spare_reg_activation_9_23), .weight_in(spare_reg_weight_8_24), .partial_sum_in(spare_reg_psum_8_24), .reg_activation(spare_reg_activation_9_24), .reg_weight(spare_reg_weight_9_24), .reg_partial_sum(spare_reg_psum_9_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_25( .activation_in(spare_reg_activation_9_24), .weight_in(spare_reg_weight_8_25), .partial_sum_in(spare_reg_psum_8_25), .reg_activation(spare_reg_activation_9_25), .reg_weight(spare_reg_weight_9_25), .reg_partial_sum(spare_reg_psum_9_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_26( .activation_in(spare_reg_activation_9_25), .weight_in(spare_reg_weight_8_26), .partial_sum_in(spare_reg_psum_8_26), .reg_activation(spare_reg_activation_9_26), .reg_weight(spare_reg_weight_9_26), .reg_partial_sum(spare_reg_psum_9_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_27( .activation_in(spare_reg_activation_9_26), .weight_in(spare_reg_weight_8_27), .partial_sum_in(spare_reg_psum_8_27), .reg_activation(spare_reg_activation_9_27), .reg_weight(spare_reg_weight_9_27), .reg_partial_sum(spare_reg_psum_9_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_28( .activation_in(spare_reg_activation_9_27), .weight_in(spare_reg_weight_8_28), .partial_sum_in(spare_reg_psum_8_28), .reg_activation(spare_reg_activation_9_28), .reg_weight(spare_reg_weight_9_28), .reg_partial_sum(spare_reg_psum_9_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_29( .activation_in(spare_reg_activation_9_28), .weight_in(spare_reg_weight_8_29), .partial_sum_in(spare_reg_psum_8_29), .reg_activation(spare_reg_activation_9_29), .reg_weight(spare_reg_weight_9_29), .reg_partial_sum(spare_reg_psum_9_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_30( .activation_in(spare_reg_activation_9_29), .weight_in(spare_reg_weight_8_30), .partial_sum_in(spare_reg_psum_8_30), .reg_activation(spare_reg_activation_9_30), .reg_weight(spare_reg_weight_9_30), .reg_partial_sum(spare_reg_psum_9_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X9_31( .activation_in(spare_reg_activation_9_30), .weight_in(spare_reg_weight_8_31), .partial_sum_in(spare_reg_psum_8_31), .reg_weight(spare_reg_weight_9_31), .reg_partial_sum(spare_reg_psum_9_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_0( .activation_in(in_activation_10), .weight_in(spare_reg_weight_9_0), .partial_sum_in(spare_reg_psum_9_0), .reg_activation(spare_reg_activation_10_0), .reg_weight(spare_reg_weight_10_0), .reg_partial_sum(spare_reg_psum_10_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_1( .activation_in(spare_reg_activation_10_0), .weight_in(spare_reg_weight_9_1), .partial_sum_in(spare_reg_psum_9_1), .reg_activation(spare_reg_activation_10_1), .reg_weight(spare_reg_weight_10_1), .reg_partial_sum(spare_reg_psum_10_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_2( .activation_in(spare_reg_activation_10_1), .weight_in(spare_reg_weight_9_2), .partial_sum_in(spare_reg_psum_9_2), .reg_activation(spare_reg_activation_10_2), .reg_weight(spare_reg_weight_10_2), .reg_partial_sum(spare_reg_psum_10_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_3( .activation_in(spare_reg_activation_10_2), .weight_in(spare_reg_weight_9_3), .partial_sum_in(spare_reg_psum_9_3), .reg_activation(spare_reg_activation_10_3), .reg_weight(spare_reg_weight_10_3), .reg_partial_sum(spare_reg_psum_10_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_4( .activation_in(spare_reg_activation_10_3), .weight_in(spare_reg_weight_9_4), .partial_sum_in(spare_reg_psum_9_4), .reg_activation(spare_reg_activation_10_4), .reg_weight(spare_reg_weight_10_4), .reg_partial_sum(spare_reg_psum_10_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_5( .activation_in(spare_reg_activation_10_4), .weight_in(spare_reg_weight_9_5), .partial_sum_in(spare_reg_psum_9_5), .reg_activation(spare_reg_activation_10_5), .reg_weight(spare_reg_weight_10_5), .reg_partial_sum(spare_reg_psum_10_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_6( .activation_in(spare_reg_activation_10_5), .weight_in(spare_reg_weight_9_6), .partial_sum_in(spare_reg_psum_9_6), .reg_activation(spare_reg_activation_10_6), .reg_weight(spare_reg_weight_10_6), .reg_partial_sum(spare_reg_psum_10_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_7( .activation_in(spare_reg_activation_10_6), .weight_in(spare_reg_weight_9_7), .partial_sum_in(spare_reg_psum_9_7), .reg_activation(spare_reg_activation_10_7), .reg_weight(spare_reg_weight_10_7), .reg_partial_sum(spare_reg_psum_10_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_8( .activation_in(spare_reg_activation_10_7), .weight_in(spare_reg_weight_9_8), .partial_sum_in(spare_reg_psum_9_8), .reg_activation(spare_reg_activation_10_8), .reg_weight(spare_reg_weight_10_8), .reg_partial_sum(spare_reg_psum_10_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_9( .activation_in(spare_reg_activation_10_8), .weight_in(spare_reg_weight_9_9), .partial_sum_in(spare_reg_psum_9_9), .reg_activation(spare_reg_activation_10_9), .reg_weight(spare_reg_weight_10_9), .reg_partial_sum(spare_reg_psum_10_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_10( .activation_in(spare_reg_activation_10_9), .weight_in(spare_reg_weight_9_10), .partial_sum_in(spare_reg_psum_9_10), .reg_activation(spare_reg_activation_10_10), .reg_weight(spare_reg_weight_10_10), .reg_partial_sum(spare_reg_psum_10_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_11( .activation_in(spare_reg_activation_10_10), .weight_in(spare_reg_weight_9_11), .partial_sum_in(spare_reg_psum_9_11), .reg_activation(spare_reg_activation_10_11), .reg_weight(spare_reg_weight_10_11), .reg_partial_sum(spare_reg_psum_10_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_12( .activation_in(spare_reg_activation_10_11), .weight_in(spare_reg_weight_9_12), .partial_sum_in(spare_reg_psum_9_12), .reg_activation(spare_reg_activation_10_12), .reg_weight(spare_reg_weight_10_12), .reg_partial_sum(spare_reg_psum_10_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_13( .activation_in(spare_reg_activation_10_12), .weight_in(spare_reg_weight_9_13), .partial_sum_in(spare_reg_psum_9_13), .reg_activation(spare_reg_activation_10_13), .reg_weight(spare_reg_weight_10_13), .reg_partial_sum(spare_reg_psum_10_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_14( .activation_in(spare_reg_activation_10_13), .weight_in(spare_reg_weight_9_14), .partial_sum_in(spare_reg_psum_9_14), .reg_activation(spare_reg_activation_10_14), .reg_weight(spare_reg_weight_10_14), .reg_partial_sum(spare_reg_psum_10_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_15( .activation_in(spare_reg_activation_10_14), .weight_in(spare_reg_weight_9_15), .partial_sum_in(spare_reg_psum_9_15), .reg_activation(spare_reg_activation_10_15), .reg_weight(spare_reg_weight_10_15), .reg_partial_sum(spare_reg_psum_10_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_16( .activation_in(spare_reg_activation_10_15), .weight_in(spare_reg_weight_9_16), .partial_sum_in(spare_reg_psum_9_16), .reg_activation(spare_reg_activation_10_16), .reg_weight(spare_reg_weight_10_16), .reg_partial_sum(spare_reg_psum_10_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_17( .activation_in(spare_reg_activation_10_16), .weight_in(spare_reg_weight_9_17), .partial_sum_in(spare_reg_psum_9_17), .reg_activation(spare_reg_activation_10_17), .reg_weight(spare_reg_weight_10_17), .reg_partial_sum(spare_reg_psum_10_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_18( .activation_in(spare_reg_activation_10_17), .weight_in(spare_reg_weight_9_18), .partial_sum_in(spare_reg_psum_9_18), .reg_activation(spare_reg_activation_10_18), .reg_weight(spare_reg_weight_10_18), .reg_partial_sum(spare_reg_psum_10_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_19( .activation_in(spare_reg_activation_10_18), .weight_in(spare_reg_weight_9_19), .partial_sum_in(spare_reg_psum_9_19), .reg_activation(spare_reg_activation_10_19), .reg_weight(spare_reg_weight_10_19), .reg_partial_sum(spare_reg_psum_10_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_20( .activation_in(spare_reg_activation_10_19), .weight_in(spare_reg_weight_9_20), .partial_sum_in(spare_reg_psum_9_20), .reg_activation(spare_reg_activation_10_20), .reg_weight(spare_reg_weight_10_20), .reg_partial_sum(spare_reg_psum_10_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_21( .activation_in(spare_reg_activation_10_20), .weight_in(spare_reg_weight_9_21), .partial_sum_in(spare_reg_psum_9_21), .reg_activation(spare_reg_activation_10_21), .reg_weight(spare_reg_weight_10_21), .reg_partial_sum(spare_reg_psum_10_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_22( .activation_in(spare_reg_activation_10_21), .weight_in(spare_reg_weight_9_22), .partial_sum_in(spare_reg_psum_9_22), .reg_activation(spare_reg_activation_10_22), .reg_weight(spare_reg_weight_10_22), .reg_partial_sum(spare_reg_psum_10_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_23( .activation_in(spare_reg_activation_10_22), .weight_in(spare_reg_weight_9_23), .partial_sum_in(spare_reg_psum_9_23), .reg_activation(spare_reg_activation_10_23), .reg_weight(spare_reg_weight_10_23), .reg_partial_sum(spare_reg_psum_10_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_24( .activation_in(spare_reg_activation_10_23), .weight_in(spare_reg_weight_9_24), .partial_sum_in(spare_reg_psum_9_24), .reg_activation(spare_reg_activation_10_24), .reg_weight(spare_reg_weight_10_24), .reg_partial_sum(spare_reg_psum_10_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_25( .activation_in(spare_reg_activation_10_24), .weight_in(spare_reg_weight_9_25), .partial_sum_in(spare_reg_psum_9_25), .reg_activation(spare_reg_activation_10_25), .reg_weight(spare_reg_weight_10_25), .reg_partial_sum(spare_reg_psum_10_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_26( .activation_in(spare_reg_activation_10_25), .weight_in(spare_reg_weight_9_26), .partial_sum_in(spare_reg_psum_9_26), .reg_activation(spare_reg_activation_10_26), .reg_weight(spare_reg_weight_10_26), .reg_partial_sum(spare_reg_psum_10_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_27( .activation_in(spare_reg_activation_10_26), .weight_in(spare_reg_weight_9_27), .partial_sum_in(spare_reg_psum_9_27), .reg_activation(spare_reg_activation_10_27), .reg_weight(spare_reg_weight_10_27), .reg_partial_sum(spare_reg_psum_10_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_28( .activation_in(spare_reg_activation_10_27), .weight_in(spare_reg_weight_9_28), .partial_sum_in(spare_reg_psum_9_28), .reg_activation(spare_reg_activation_10_28), .reg_weight(spare_reg_weight_10_28), .reg_partial_sum(spare_reg_psum_10_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_29( .activation_in(spare_reg_activation_10_28), .weight_in(spare_reg_weight_9_29), .partial_sum_in(spare_reg_psum_9_29), .reg_activation(spare_reg_activation_10_29), .reg_weight(spare_reg_weight_10_29), .reg_partial_sum(spare_reg_psum_10_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_30( .activation_in(spare_reg_activation_10_29), .weight_in(spare_reg_weight_9_30), .partial_sum_in(spare_reg_psum_9_30), .reg_activation(spare_reg_activation_10_30), .reg_weight(spare_reg_weight_10_30), .reg_partial_sum(spare_reg_psum_10_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X10_31( .activation_in(spare_reg_activation_10_30), .weight_in(spare_reg_weight_9_31), .partial_sum_in(spare_reg_psum_9_31), .reg_weight(spare_reg_weight_10_31), .reg_partial_sum(spare_reg_psum_10_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_0( .activation_in(in_activation_11), .weight_in(spare_reg_weight_10_0), .partial_sum_in(spare_reg_psum_10_0), .reg_activation(spare_reg_activation_11_0), .reg_weight(spare_reg_weight_11_0), .reg_partial_sum(spare_reg_psum_11_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_1( .activation_in(spare_reg_activation_11_0), .weight_in(spare_reg_weight_10_1), .partial_sum_in(spare_reg_psum_10_1), .reg_activation(spare_reg_activation_11_1), .reg_weight(spare_reg_weight_11_1), .reg_partial_sum(spare_reg_psum_11_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_2( .activation_in(spare_reg_activation_11_1), .weight_in(spare_reg_weight_10_2), .partial_sum_in(spare_reg_psum_10_2), .reg_activation(spare_reg_activation_11_2), .reg_weight(spare_reg_weight_11_2), .reg_partial_sum(spare_reg_psum_11_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_3( .activation_in(spare_reg_activation_11_2), .weight_in(spare_reg_weight_10_3), .partial_sum_in(spare_reg_psum_10_3), .reg_activation(spare_reg_activation_11_3), .reg_weight(spare_reg_weight_11_3), .reg_partial_sum(spare_reg_psum_11_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_4( .activation_in(spare_reg_activation_11_3), .weight_in(spare_reg_weight_10_4), .partial_sum_in(spare_reg_psum_10_4), .reg_activation(spare_reg_activation_11_4), .reg_weight(spare_reg_weight_11_4), .reg_partial_sum(spare_reg_psum_11_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_5( .activation_in(spare_reg_activation_11_4), .weight_in(spare_reg_weight_10_5), .partial_sum_in(spare_reg_psum_10_5), .reg_activation(spare_reg_activation_11_5), .reg_weight(spare_reg_weight_11_5), .reg_partial_sum(spare_reg_psum_11_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_6( .activation_in(spare_reg_activation_11_5), .weight_in(spare_reg_weight_10_6), .partial_sum_in(spare_reg_psum_10_6), .reg_activation(spare_reg_activation_11_6), .reg_weight(spare_reg_weight_11_6), .reg_partial_sum(spare_reg_psum_11_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_7( .activation_in(spare_reg_activation_11_6), .weight_in(spare_reg_weight_10_7), .partial_sum_in(spare_reg_psum_10_7), .reg_activation(spare_reg_activation_11_7), .reg_weight(spare_reg_weight_11_7), .reg_partial_sum(spare_reg_psum_11_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_8( .activation_in(spare_reg_activation_11_7), .weight_in(spare_reg_weight_10_8), .partial_sum_in(spare_reg_psum_10_8), .reg_activation(spare_reg_activation_11_8), .reg_weight(spare_reg_weight_11_8), .reg_partial_sum(spare_reg_psum_11_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_9( .activation_in(spare_reg_activation_11_8), .weight_in(spare_reg_weight_10_9), .partial_sum_in(spare_reg_psum_10_9), .reg_activation(spare_reg_activation_11_9), .reg_weight(spare_reg_weight_11_9), .reg_partial_sum(spare_reg_psum_11_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_10( .activation_in(spare_reg_activation_11_9), .weight_in(spare_reg_weight_10_10), .partial_sum_in(spare_reg_psum_10_10), .reg_activation(spare_reg_activation_11_10), .reg_weight(spare_reg_weight_11_10), .reg_partial_sum(spare_reg_psum_11_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_11( .activation_in(spare_reg_activation_11_10), .weight_in(spare_reg_weight_10_11), .partial_sum_in(spare_reg_psum_10_11), .reg_activation(spare_reg_activation_11_11), .reg_weight(spare_reg_weight_11_11), .reg_partial_sum(spare_reg_psum_11_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_12( .activation_in(spare_reg_activation_11_11), .weight_in(spare_reg_weight_10_12), .partial_sum_in(spare_reg_psum_10_12), .reg_activation(spare_reg_activation_11_12), .reg_weight(spare_reg_weight_11_12), .reg_partial_sum(spare_reg_psum_11_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_13( .activation_in(spare_reg_activation_11_12), .weight_in(spare_reg_weight_10_13), .partial_sum_in(spare_reg_psum_10_13), .reg_activation(spare_reg_activation_11_13), .reg_weight(spare_reg_weight_11_13), .reg_partial_sum(spare_reg_psum_11_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_14( .activation_in(spare_reg_activation_11_13), .weight_in(spare_reg_weight_10_14), .partial_sum_in(spare_reg_psum_10_14), .reg_activation(spare_reg_activation_11_14), .reg_weight(spare_reg_weight_11_14), .reg_partial_sum(spare_reg_psum_11_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_15( .activation_in(spare_reg_activation_11_14), .weight_in(spare_reg_weight_10_15), .partial_sum_in(spare_reg_psum_10_15), .reg_activation(spare_reg_activation_11_15), .reg_weight(spare_reg_weight_11_15), .reg_partial_sum(spare_reg_psum_11_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_16( .activation_in(spare_reg_activation_11_15), .weight_in(spare_reg_weight_10_16), .partial_sum_in(spare_reg_psum_10_16), .reg_activation(spare_reg_activation_11_16), .reg_weight(spare_reg_weight_11_16), .reg_partial_sum(spare_reg_psum_11_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_17( .activation_in(spare_reg_activation_11_16), .weight_in(spare_reg_weight_10_17), .partial_sum_in(spare_reg_psum_10_17), .reg_activation(spare_reg_activation_11_17), .reg_weight(spare_reg_weight_11_17), .reg_partial_sum(spare_reg_psum_11_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_18( .activation_in(spare_reg_activation_11_17), .weight_in(spare_reg_weight_10_18), .partial_sum_in(spare_reg_psum_10_18), .reg_activation(spare_reg_activation_11_18), .reg_weight(spare_reg_weight_11_18), .reg_partial_sum(spare_reg_psum_11_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_19( .activation_in(spare_reg_activation_11_18), .weight_in(spare_reg_weight_10_19), .partial_sum_in(spare_reg_psum_10_19), .reg_activation(spare_reg_activation_11_19), .reg_weight(spare_reg_weight_11_19), .reg_partial_sum(spare_reg_psum_11_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_20( .activation_in(spare_reg_activation_11_19), .weight_in(spare_reg_weight_10_20), .partial_sum_in(spare_reg_psum_10_20), .reg_activation(spare_reg_activation_11_20), .reg_weight(spare_reg_weight_11_20), .reg_partial_sum(spare_reg_psum_11_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_21( .activation_in(spare_reg_activation_11_20), .weight_in(spare_reg_weight_10_21), .partial_sum_in(spare_reg_psum_10_21), .reg_activation(spare_reg_activation_11_21), .reg_weight(spare_reg_weight_11_21), .reg_partial_sum(spare_reg_psum_11_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_22( .activation_in(spare_reg_activation_11_21), .weight_in(spare_reg_weight_10_22), .partial_sum_in(spare_reg_psum_10_22), .reg_activation(spare_reg_activation_11_22), .reg_weight(spare_reg_weight_11_22), .reg_partial_sum(spare_reg_psum_11_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_23( .activation_in(spare_reg_activation_11_22), .weight_in(spare_reg_weight_10_23), .partial_sum_in(spare_reg_psum_10_23), .reg_activation(spare_reg_activation_11_23), .reg_weight(spare_reg_weight_11_23), .reg_partial_sum(spare_reg_psum_11_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_24( .activation_in(spare_reg_activation_11_23), .weight_in(spare_reg_weight_10_24), .partial_sum_in(spare_reg_psum_10_24), .reg_activation(spare_reg_activation_11_24), .reg_weight(spare_reg_weight_11_24), .reg_partial_sum(spare_reg_psum_11_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_25( .activation_in(spare_reg_activation_11_24), .weight_in(spare_reg_weight_10_25), .partial_sum_in(spare_reg_psum_10_25), .reg_activation(spare_reg_activation_11_25), .reg_weight(spare_reg_weight_11_25), .reg_partial_sum(spare_reg_psum_11_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_26( .activation_in(spare_reg_activation_11_25), .weight_in(spare_reg_weight_10_26), .partial_sum_in(spare_reg_psum_10_26), .reg_activation(spare_reg_activation_11_26), .reg_weight(spare_reg_weight_11_26), .reg_partial_sum(spare_reg_psum_11_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_27( .activation_in(spare_reg_activation_11_26), .weight_in(spare_reg_weight_10_27), .partial_sum_in(spare_reg_psum_10_27), .reg_activation(spare_reg_activation_11_27), .reg_weight(spare_reg_weight_11_27), .reg_partial_sum(spare_reg_psum_11_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_28( .activation_in(spare_reg_activation_11_27), .weight_in(spare_reg_weight_10_28), .partial_sum_in(spare_reg_psum_10_28), .reg_activation(spare_reg_activation_11_28), .reg_weight(spare_reg_weight_11_28), .reg_partial_sum(spare_reg_psum_11_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_29( .activation_in(spare_reg_activation_11_28), .weight_in(spare_reg_weight_10_29), .partial_sum_in(spare_reg_psum_10_29), .reg_activation(spare_reg_activation_11_29), .reg_weight(spare_reg_weight_11_29), .reg_partial_sum(spare_reg_psum_11_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_30( .activation_in(spare_reg_activation_11_29), .weight_in(spare_reg_weight_10_30), .partial_sum_in(spare_reg_psum_10_30), .reg_activation(spare_reg_activation_11_30), .reg_weight(spare_reg_weight_11_30), .reg_partial_sum(spare_reg_psum_11_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X11_31( .activation_in(spare_reg_activation_11_30), .weight_in(spare_reg_weight_10_31), .partial_sum_in(spare_reg_psum_10_31), .reg_weight(spare_reg_weight_11_31), .reg_partial_sum(spare_reg_psum_11_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_0( .activation_in(in_activation_12), .weight_in(spare_reg_weight_11_0), .partial_sum_in(spare_reg_psum_11_0), .reg_activation(spare_reg_activation_12_0), .reg_weight(spare_reg_weight_12_0), .reg_partial_sum(spare_reg_psum_12_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_1( .activation_in(spare_reg_activation_12_0), .weight_in(spare_reg_weight_11_1), .partial_sum_in(spare_reg_psum_11_1), .reg_activation(spare_reg_activation_12_1), .reg_weight(spare_reg_weight_12_1), .reg_partial_sum(spare_reg_psum_12_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_2( .activation_in(spare_reg_activation_12_1), .weight_in(spare_reg_weight_11_2), .partial_sum_in(spare_reg_psum_11_2), .reg_activation(spare_reg_activation_12_2), .reg_weight(spare_reg_weight_12_2), .reg_partial_sum(spare_reg_psum_12_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_3( .activation_in(spare_reg_activation_12_2), .weight_in(spare_reg_weight_11_3), .partial_sum_in(spare_reg_psum_11_3), .reg_activation(spare_reg_activation_12_3), .reg_weight(spare_reg_weight_12_3), .reg_partial_sum(spare_reg_psum_12_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_4( .activation_in(spare_reg_activation_12_3), .weight_in(spare_reg_weight_11_4), .partial_sum_in(spare_reg_psum_11_4), .reg_activation(spare_reg_activation_12_4), .reg_weight(spare_reg_weight_12_4), .reg_partial_sum(spare_reg_psum_12_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_5( .activation_in(spare_reg_activation_12_4), .weight_in(spare_reg_weight_11_5), .partial_sum_in(spare_reg_psum_11_5), .reg_activation(spare_reg_activation_12_5), .reg_weight(spare_reg_weight_12_5), .reg_partial_sum(spare_reg_psum_12_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_6( .activation_in(spare_reg_activation_12_5), .weight_in(spare_reg_weight_11_6), .partial_sum_in(spare_reg_psum_11_6), .reg_activation(spare_reg_activation_12_6), .reg_weight(spare_reg_weight_12_6), .reg_partial_sum(spare_reg_psum_12_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_7( .activation_in(spare_reg_activation_12_6), .weight_in(spare_reg_weight_11_7), .partial_sum_in(spare_reg_psum_11_7), .reg_activation(spare_reg_activation_12_7), .reg_weight(spare_reg_weight_12_7), .reg_partial_sum(spare_reg_psum_12_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_8( .activation_in(spare_reg_activation_12_7), .weight_in(spare_reg_weight_11_8), .partial_sum_in(spare_reg_psum_11_8), .reg_activation(spare_reg_activation_12_8), .reg_weight(spare_reg_weight_12_8), .reg_partial_sum(spare_reg_psum_12_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_9( .activation_in(spare_reg_activation_12_8), .weight_in(spare_reg_weight_11_9), .partial_sum_in(spare_reg_psum_11_9), .reg_activation(spare_reg_activation_12_9), .reg_weight(spare_reg_weight_12_9), .reg_partial_sum(spare_reg_psum_12_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_10( .activation_in(spare_reg_activation_12_9), .weight_in(spare_reg_weight_11_10), .partial_sum_in(spare_reg_psum_11_10), .reg_activation(spare_reg_activation_12_10), .reg_weight(spare_reg_weight_12_10), .reg_partial_sum(spare_reg_psum_12_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_11( .activation_in(spare_reg_activation_12_10), .weight_in(spare_reg_weight_11_11), .partial_sum_in(spare_reg_psum_11_11), .reg_activation(spare_reg_activation_12_11), .reg_weight(spare_reg_weight_12_11), .reg_partial_sum(spare_reg_psum_12_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_12( .activation_in(spare_reg_activation_12_11), .weight_in(spare_reg_weight_11_12), .partial_sum_in(spare_reg_psum_11_12), .reg_activation(spare_reg_activation_12_12), .reg_weight(spare_reg_weight_12_12), .reg_partial_sum(spare_reg_psum_12_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_13( .activation_in(spare_reg_activation_12_12), .weight_in(spare_reg_weight_11_13), .partial_sum_in(spare_reg_psum_11_13), .reg_activation(spare_reg_activation_12_13), .reg_weight(spare_reg_weight_12_13), .reg_partial_sum(spare_reg_psum_12_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_14( .activation_in(spare_reg_activation_12_13), .weight_in(spare_reg_weight_11_14), .partial_sum_in(spare_reg_psum_11_14), .reg_activation(spare_reg_activation_12_14), .reg_weight(spare_reg_weight_12_14), .reg_partial_sum(spare_reg_psum_12_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_15( .activation_in(spare_reg_activation_12_14), .weight_in(spare_reg_weight_11_15), .partial_sum_in(spare_reg_psum_11_15), .reg_activation(spare_reg_activation_12_15), .reg_weight(spare_reg_weight_12_15), .reg_partial_sum(spare_reg_psum_12_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_16( .activation_in(spare_reg_activation_12_15), .weight_in(spare_reg_weight_11_16), .partial_sum_in(spare_reg_psum_11_16), .reg_activation(spare_reg_activation_12_16), .reg_weight(spare_reg_weight_12_16), .reg_partial_sum(spare_reg_psum_12_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_17( .activation_in(spare_reg_activation_12_16), .weight_in(spare_reg_weight_11_17), .partial_sum_in(spare_reg_psum_11_17), .reg_activation(spare_reg_activation_12_17), .reg_weight(spare_reg_weight_12_17), .reg_partial_sum(spare_reg_psum_12_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_18( .activation_in(spare_reg_activation_12_17), .weight_in(spare_reg_weight_11_18), .partial_sum_in(spare_reg_psum_11_18), .reg_activation(spare_reg_activation_12_18), .reg_weight(spare_reg_weight_12_18), .reg_partial_sum(spare_reg_psum_12_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_19( .activation_in(spare_reg_activation_12_18), .weight_in(spare_reg_weight_11_19), .partial_sum_in(spare_reg_psum_11_19), .reg_activation(spare_reg_activation_12_19), .reg_weight(spare_reg_weight_12_19), .reg_partial_sum(spare_reg_psum_12_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_20( .activation_in(spare_reg_activation_12_19), .weight_in(spare_reg_weight_11_20), .partial_sum_in(spare_reg_psum_11_20), .reg_activation(spare_reg_activation_12_20), .reg_weight(spare_reg_weight_12_20), .reg_partial_sum(spare_reg_psum_12_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_21( .activation_in(spare_reg_activation_12_20), .weight_in(spare_reg_weight_11_21), .partial_sum_in(spare_reg_psum_11_21), .reg_activation(spare_reg_activation_12_21), .reg_weight(spare_reg_weight_12_21), .reg_partial_sum(spare_reg_psum_12_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_22( .activation_in(spare_reg_activation_12_21), .weight_in(spare_reg_weight_11_22), .partial_sum_in(spare_reg_psum_11_22), .reg_activation(spare_reg_activation_12_22), .reg_weight(spare_reg_weight_12_22), .reg_partial_sum(spare_reg_psum_12_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_23( .activation_in(spare_reg_activation_12_22), .weight_in(spare_reg_weight_11_23), .partial_sum_in(spare_reg_psum_11_23), .reg_activation(spare_reg_activation_12_23), .reg_weight(spare_reg_weight_12_23), .reg_partial_sum(spare_reg_psum_12_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_24( .activation_in(spare_reg_activation_12_23), .weight_in(spare_reg_weight_11_24), .partial_sum_in(spare_reg_psum_11_24), .reg_activation(spare_reg_activation_12_24), .reg_weight(spare_reg_weight_12_24), .reg_partial_sum(spare_reg_psum_12_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_25( .activation_in(spare_reg_activation_12_24), .weight_in(spare_reg_weight_11_25), .partial_sum_in(spare_reg_psum_11_25), .reg_activation(spare_reg_activation_12_25), .reg_weight(spare_reg_weight_12_25), .reg_partial_sum(spare_reg_psum_12_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_26( .activation_in(spare_reg_activation_12_25), .weight_in(spare_reg_weight_11_26), .partial_sum_in(spare_reg_psum_11_26), .reg_activation(spare_reg_activation_12_26), .reg_weight(spare_reg_weight_12_26), .reg_partial_sum(spare_reg_psum_12_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_27( .activation_in(spare_reg_activation_12_26), .weight_in(spare_reg_weight_11_27), .partial_sum_in(spare_reg_psum_11_27), .reg_activation(spare_reg_activation_12_27), .reg_weight(spare_reg_weight_12_27), .reg_partial_sum(spare_reg_psum_12_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_28( .activation_in(spare_reg_activation_12_27), .weight_in(spare_reg_weight_11_28), .partial_sum_in(spare_reg_psum_11_28), .reg_activation(spare_reg_activation_12_28), .reg_weight(spare_reg_weight_12_28), .reg_partial_sum(spare_reg_psum_12_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_29( .activation_in(spare_reg_activation_12_28), .weight_in(spare_reg_weight_11_29), .partial_sum_in(spare_reg_psum_11_29), .reg_activation(spare_reg_activation_12_29), .reg_weight(spare_reg_weight_12_29), .reg_partial_sum(spare_reg_psum_12_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_30( .activation_in(spare_reg_activation_12_29), .weight_in(spare_reg_weight_11_30), .partial_sum_in(spare_reg_psum_11_30), .reg_activation(spare_reg_activation_12_30), .reg_weight(spare_reg_weight_12_30), .reg_partial_sum(spare_reg_psum_12_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X12_31( .activation_in(spare_reg_activation_12_30), .weight_in(spare_reg_weight_11_31), .partial_sum_in(spare_reg_psum_11_31), .reg_weight(spare_reg_weight_12_31), .reg_partial_sum(spare_reg_psum_12_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_0( .activation_in(in_activation_13), .weight_in(spare_reg_weight_12_0), .partial_sum_in(spare_reg_psum_12_0), .reg_activation(spare_reg_activation_13_0), .reg_weight(spare_reg_weight_13_0), .reg_partial_sum(spare_reg_psum_13_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_1( .activation_in(spare_reg_activation_13_0), .weight_in(spare_reg_weight_12_1), .partial_sum_in(spare_reg_psum_12_1), .reg_activation(spare_reg_activation_13_1), .reg_weight(spare_reg_weight_13_1), .reg_partial_sum(spare_reg_psum_13_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_2( .activation_in(spare_reg_activation_13_1), .weight_in(spare_reg_weight_12_2), .partial_sum_in(spare_reg_psum_12_2), .reg_activation(spare_reg_activation_13_2), .reg_weight(spare_reg_weight_13_2), .reg_partial_sum(spare_reg_psum_13_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_3( .activation_in(spare_reg_activation_13_2), .weight_in(spare_reg_weight_12_3), .partial_sum_in(spare_reg_psum_12_3), .reg_activation(spare_reg_activation_13_3), .reg_weight(spare_reg_weight_13_3), .reg_partial_sum(spare_reg_psum_13_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_4( .activation_in(spare_reg_activation_13_3), .weight_in(spare_reg_weight_12_4), .partial_sum_in(spare_reg_psum_12_4), .reg_activation(spare_reg_activation_13_4), .reg_weight(spare_reg_weight_13_4), .reg_partial_sum(spare_reg_psum_13_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_5( .activation_in(spare_reg_activation_13_4), .weight_in(spare_reg_weight_12_5), .partial_sum_in(spare_reg_psum_12_5), .reg_activation(spare_reg_activation_13_5), .reg_weight(spare_reg_weight_13_5), .reg_partial_sum(spare_reg_psum_13_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_6( .activation_in(spare_reg_activation_13_5), .weight_in(spare_reg_weight_12_6), .partial_sum_in(spare_reg_psum_12_6), .reg_activation(spare_reg_activation_13_6), .reg_weight(spare_reg_weight_13_6), .reg_partial_sum(spare_reg_psum_13_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_7( .activation_in(spare_reg_activation_13_6), .weight_in(spare_reg_weight_12_7), .partial_sum_in(spare_reg_psum_12_7), .reg_activation(spare_reg_activation_13_7), .reg_weight(spare_reg_weight_13_7), .reg_partial_sum(spare_reg_psum_13_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_8( .activation_in(spare_reg_activation_13_7), .weight_in(spare_reg_weight_12_8), .partial_sum_in(spare_reg_psum_12_8), .reg_activation(spare_reg_activation_13_8), .reg_weight(spare_reg_weight_13_8), .reg_partial_sum(spare_reg_psum_13_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_9( .activation_in(spare_reg_activation_13_8), .weight_in(spare_reg_weight_12_9), .partial_sum_in(spare_reg_psum_12_9), .reg_activation(spare_reg_activation_13_9), .reg_weight(spare_reg_weight_13_9), .reg_partial_sum(spare_reg_psum_13_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_10( .activation_in(spare_reg_activation_13_9), .weight_in(spare_reg_weight_12_10), .partial_sum_in(spare_reg_psum_12_10), .reg_activation(spare_reg_activation_13_10), .reg_weight(spare_reg_weight_13_10), .reg_partial_sum(spare_reg_psum_13_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_11( .activation_in(spare_reg_activation_13_10), .weight_in(spare_reg_weight_12_11), .partial_sum_in(spare_reg_psum_12_11), .reg_activation(spare_reg_activation_13_11), .reg_weight(spare_reg_weight_13_11), .reg_partial_sum(spare_reg_psum_13_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_12( .activation_in(spare_reg_activation_13_11), .weight_in(spare_reg_weight_12_12), .partial_sum_in(spare_reg_psum_12_12), .reg_activation(spare_reg_activation_13_12), .reg_weight(spare_reg_weight_13_12), .reg_partial_sum(spare_reg_psum_13_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_13( .activation_in(spare_reg_activation_13_12), .weight_in(spare_reg_weight_12_13), .partial_sum_in(spare_reg_psum_12_13), .reg_activation(spare_reg_activation_13_13), .reg_weight(spare_reg_weight_13_13), .reg_partial_sum(spare_reg_psum_13_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_14( .activation_in(spare_reg_activation_13_13), .weight_in(spare_reg_weight_12_14), .partial_sum_in(spare_reg_psum_12_14), .reg_activation(spare_reg_activation_13_14), .reg_weight(spare_reg_weight_13_14), .reg_partial_sum(spare_reg_psum_13_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_15( .activation_in(spare_reg_activation_13_14), .weight_in(spare_reg_weight_12_15), .partial_sum_in(spare_reg_psum_12_15), .reg_activation(spare_reg_activation_13_15), .reg_weight(spare_reg_weight_13_15), .reg_partial_sum(spare_reg_psum_13_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_16( .activation_in(spare_reg_activation_13_15), .weight_in(spare_reg_weight_12_16), .partial_sum_in(spare_reg_psum_12_16), .reg_activation(spare_reg_activation_13_16), .reg_weight(spare_reg_weight_13_16), .reg_partial_sum(spare_reg_psum_13_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_17( .activation_in(spare_reg_activation_13_16), .weight_in(spare_reg_weight_12_17), .partial_sum_in(spare_reg_psum_12_17), .reg_activation(spare_reg_activation_13_17), .reg_weight(spare_reg_weight_13_17), .reg_partial_sum(spare_reg_psum_13_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_18( .activation_in(spare_reg_activation_13_17), .weight_in(spare_reg_weight_12_18), .partial_sum_in(spare_reg_psum_12_18), .reg_activation(spare_reg_activation_13_18), .reg_weight(spare_reg_weight_13_18), .reg_partial_sum(spare_reg_psum_13_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_19( .activation_in(spare_reg_activation_13_18), .weight_in(spare_reg_weight_12_19), .partial_sum_in(spare_reg_psum_12_19), .reg_activation(spare_reg_activation_13_19), .reg_weight(spare_reg_weight_13_19), .reg_partial_sum(spare_reg_psum_13_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_20( .activation_in(spare_reg_activation_13_19), .weight_in(spare_reg_weight_12_20), .partial_sum_in(spare_reg_psum_12_20), .reg_activation(spare_reg_activation_13_20), .reg_weight(spare_reg_weight_13_20), .reg_partial_sum(spare_reg_psum_13_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_21( .activation_in(spare_reg_activation_13_20), .weight_in(spare_reg_weight_12_21), .partial_sum_in(spare_reg_psum_12_21), .reg_activation(spare_reg_activation_13_21), .reg_weight(spare_reg_weight_13_21), .reg_partial_sum(spare_reg_psum_13_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_22( .activation_in(spare_reg_activation_13_21), .weight_in(spare_reg_weight_12_22), .partial_sum_in(spare_reg_psum_12_22), .reg_activation(spare_reg_activation_13_22), .reg_weight(spare_reg_weight_13_22), .reg_partial_sum(spare_reg_psum_13_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_23( .activation_in(spare_reg_activation_13_22), .weight_in(spare_reg_weight_12_23), .partial_sum_in(spare_reg_psum_12_23), .reg_activation(spare_reg_activation_13_23), .reg_weight(spare_reg_weight_13_23), .reg_partial_sum(spare_reg_psum_13_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_24( .activation_in(spare_reg_activation_13_23), .weight_in(spare_reg_weight_12_24), .partial_sum_in(spare_reg_psum_12_24), .reg_activation(spare_reg_activation_13_24), .reg_weight(spare_reg_weight_13_24), .reg_partial_sum(spare_reg_psum_13_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_25( .activation_in(spare_reg_activation_13_24), .weight_in(spare_reg_weight_12_25), .partial_sum_in(spare_reg_psum_12_25), .reg_activation(spare_reg_activation_13_25), .reg_weight(spare_reg_weight_13_25), .reg_partial_sum(spare_reg_psum_13_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_26( .activation_in(spare_reg_activation_13_25), .weight_in(spare_reg_weight_12_26), .partial_sum_in(spare_reg_psum_12_26), .reg_activation(spare_reg_activation_13_26), .reg_weight(spare_reg_weight_13_26), .reg_partial_sum(spare_reg_psum_13_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_27( .activation_in(spare_reg_activation_13_26), .weight_in(spare_reg_weight_12_27), .partial_sum_in(spare_reg_psum_12_27), .reg_activation(spare_reg_activation_13_27), .reg_weight(spare_reg_weight_13_27), .reg_partial_sum(spare_reg_psum_13_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_28( .activation_in(spare_reg_activation_13_27), .weight_in(spare_reg_weight_12_28), .partial_sum_in(spare_reg_psum_12_28), .reg_activation(spare_reg_activation_13_28), .reg_weight(spare_reg_weight_13_28), .reg_partial_sum(spare_reg_psum_13_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_29( .activation_in(spare_reg_activation_13_28), .weight_in(spare_reg_weight_12_29), .partial_sum_in(spare_reg_psum_12_29), .reg_activation(spare_reg_activation_13_29), .reg_weight(spare_reg_weight_13_29), .reg_partial_sum(spare_reg_psum_13_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_30( .activation_in(spare_reg_activation_13_29), .weight_in(spare_reg_weight_12_30), .partial_sum_in(spare_reg_psum_12_30), .reg_activation(spare_reg_activation_13_30), .reg_weight(spare_reg_weight_13_30), .reg_partial_sum(spare_reg_psum_13_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X13_31( .activation_in(spare_reg_activation_13_30), .weight_in(spare_reg_weight_12_31), .partial_sum_in(spare_reg_psum_12_31), .reg_weight(spare_reg_weight_13_31), .reg_partial_sum(spare_reg_psum_13_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_0( .activation_in(in_activation_14), .weight_in(spare_reg_weight_13_0), .partial_sum_in(spare_reg_psum_13_0), .reg_activation(spare_reg_activation_14_0), .reg_weight(spare_reg_weight_14_0), .reg_partial_sum(spare_reg_psum_14_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_1( .activation_in(spare_reg_activation_14_0), .weight_in(spare_reg_weight_13_1), .partial_sum_in(spare_reg_psum_13_1), .reg_activation(spare_reg_activation_14_1), .reg_weight(spare_reg_weight_14_1), .reg_partial_sum(spare_reg_psum_14_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_2( .activation_in(spare_reg_activation_14_1), .weight_in(spare_reg_weight_13_2), .partial_sum_in(spare_reg_psum_13_2), .reg_activation(spare_reg_activation_14_2), .reg_weight(spare_reg_weight_14_2), .reg_partial_sum(spare_reg_psum_14_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_3( .activation_in(spare_reg_activation_14_2), .weight_in(spare_reg_weight_13_3), .partial_sum_in(spare_reg_psum_13_3), .reg_activation(spare_reg_activation_14_3), .reg_weight(spare_reg_weight_14_3), .reg_partial_sum(spare_reg_psum_14_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_4( .activation_in(spare_reg_activation_14_3), .weight_in(spare_reg_weight_13_4), .partial_sum_in(spare_reg_psum_13_4), .reg_activation(spare_reg_activation_14_4), .reg_weight(spare_reg_weight_14_4), .reg_partial_sum(spare_reg_psum_14_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_5( .activation_in(spare_reg_activation_14_4), .weight_in(spare_reg_weight_13_5), .partial_sum_in(spare_reg_psum_13_5), .reg_activation(spare_reg_activation_14_5), .reg_weight(spare_reg_weight_14_5), .reg_partial_sum(spare_reg_psum_14_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_6( .activation_in(spare_reg_activation_14_5), .weight_in(spare_reg_weight_13_6), .partial_sum_in(spare_reg_psum_13_6), .reg_activation(spare_reg_activation_14_6), .reg_weight(spare_reg_weight_14_6), .reg_partial_sum(spare_reg_psum_14_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_7( .activation_in(spare_reg_activation_14_6), .weight_in(spare_reg_weight_13_7), .partial_sum_in(spare_reg_psum_13_7), .reg_activation(spare_reg_activation_14_7), .reg_weight(spare_reg_weight_14_7), .reg_partial_sum(spare_reg_psum_14_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_8( .activation_in(spare_reg_activation_14_7), .weight_in(spare_reg_weight_13_8), .partial_sum_in(spare_reg_psum_13_8), .reg_activation(spare_reg_activation_14_8), .reg_weight(spare_reg_weight_14_8), .reg_partial_sum(spare_reg_psum_14_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_9( .activation_in(spare_reg_activation_14_8), .weight_in(spare_reg_weight_13_9), .partial_sum_in(spare_reg_psum_13_9), .reg_activation(spare_reg_activation_14_9), .reg_weight(spare_reg_weight_14_9), .reg_partial_sum(spare_reg_psum_14_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_10( .activation_in(spare_reg_activation_14_9), .weight_in(spare_reg_weight_13_10), .partial_sum_in(spare_reg_psum_13_10), .reg_activation(spare_reg_activation_14_10), .reg_weight(spare_reg_weight_14_10), .reg_partial_sum(spare_reg_psum_14_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_11( .activation_in(spare_reg_activation_14_10), .weight_in(spare_reg_weight_13_11), .partial_sum_in(spare_reg_psum_13_11), .reg_activation(spare_reg_activation_14_11), .reg_weight(spare_reg_weight_14_11), .reg_partial_sum(spare_reg_psum_14_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_12( .activation_in(spare_reg_activation_14_11), .weight_in(spare_reg_weight_13_12), .partial_sum_in(spare_reg_psum_13_12), .reg_activation(spare_reg_activation_14_12), .reg_weight(spare_reg_weight_14_12), .reg_partial_sum(spare_reg_psum_14_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_13( .activation_in(spare_reg_activation_14_12), .weight_in(spare_reg_weight_13_13), .partial_sum_in(spare_reg_psum_13_13), .reg_activation(spare_reg_activation_14_13), .reg_weight(spare_reg_weight_14_13), .reg_partial_sum(spare_reg_psum_14_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_14( .activation_in(spare_reg_activation_14_13), .weight_in(spare_reg_weight_13_14), .partial_sum_in(spare_reg_psum_13_14), .reg_activation(spare_reg_activation_14_14), .reg_weight(spare_reg_weight_14_14), .reg_partial_sum(spare_reg_psum_14_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_15( .activation_in(spare_reg_activation_14_14), .weight_in(spare_reg_weight_13_15), .partial_sum_in(spare_reg_psum_13_15), .reg_activation(spare_reg_activation_14_15), .reg_weight(spare_reg_weight_14_15), .reg_partial_sum(spare_reg_psum_14_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_16( .activation_in(spare_reg_activation_14_15), .weight_in(spare_reg_weight_13_16), .partial_sum_in(spare_reg_psum_13_16), .reg_activation(spare_reg_activation_14_16), .reg_weight(spare_reg_weight_14_16), .reg_partial_sum(spare_reg_psum_14_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_17( .activation_in(spare_reg_activation_14_16), .weight_in(spare_reg_weight_13_17), .partial_sum_in(spare_reg_psum_13_17), .reg_activation(spare_reg_activation_14_17), .reg_weight(spare_reg_weight_14_17), .reg_partial_sum(spare_reg_psum_14_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_18( .activation_in(spare_reg_activation_14_17), .weight_in(spare_reg_weight_13_18), .partial_sum_in(spare_reg_psum_13_18), .reg_activation(spare_reg_activation_14_18), .reg_weight(spare_reg_weight_14_18), .reg_partial_sum(spare_reg_psum_14_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_19( .activation_in(spare_reg_activation_14_18), .weight_in(spare_reg_weight_13_19), .partial_sum_in(spare_reg_psum_13_19), .reg_activation(spare_reg_activation_14_19), .reg_weight(spare_reg_weight_14_19), .reg_partial_sum(spare_reg_psum_14_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_20( .activation_in(spare_reg_activation_14_19), .weight_in(spare_reg_weight_13_20), .partial_sum_in(spare_reg_psum_13_20), .reg_activation(spare_reg_activation_14_20), .reg_weight(spare_reg_weight_14_20), .reg_partial_sum(spare_reg_psum_14_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_21( .activation_in(spare_reg_activation_14_20), .weight_in(spare_reg_weight_13_21), .partial_sum_in(spare_reg_psum_13_21), .reg_activation(spare_reg_activation_14_21), .reg_weight(spare_reg_weight_14_21), .reg_partial_sum(spare_reg_psum_14_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_22( .activation_in(spare_reg_activation_14_21), .weight_in(spare_reg_weight_13_22), .partial_sum_in(spare_reg_psum_13_22), .reg_activation(spare_reg_activation_14_22), .reg_weight(spare_reg_weight_14_22), .reg_partial_sum(spare_reg_psum_14_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_23( .activation_in(spare_reg_activation_14_22), .weight_in(spare_reg_weight_13_23), .partial_sum_in(spare_reg_psum_13_23), .reg_activation(spare_reg_activation_14_23), .reg_weight(spare_reg_weight_14_23), .reg_partial_sum(spare_reg_psum_14_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_24( .activation_in(spare_reg_activation_14_23), .weight_in(spare_reg_weight_13_24), .partial_sum_in(spare_reg_psum_13_24), .reg_activation(spare_reg_activation_14_24), .reg_weight(spare_reg_weight_14_24), .reg_partial_sum(spare_reg_psum_14_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_25( .activation_in(spare_reg_activation_14_24), .weight_in(spare_reg_weight_13_25), .partial_sum_in(spare_reg_psum_13_25), .reg_activation(spare_reg_activation_14_25), .reg_weight(spare_reg_weight_14_25), .reg_partial_sum(spare_reg_psum_14_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_26( .activation_in(spare_reg_activation_14_25), .weight_in(spare_reg_weight_13_26), .partial_sum_in(spare_reg_psum_13_26), .reg_activation(spare_reg_activation_14_26), .reg_weight(spare_reg_weight_14_26), .reg_partial_sum(spare_reg_psum_14_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_27( .activation_in(spare_reg_activation_14_26), .weight_in(spare_reg_weight_13_27), .partial_sum_in(spare_reg_psum_13_27), .reg_activation(spare_reg_activation_14_27), .reg_weight(spare_reg_weight_14_27), .reg_partial_sum(spare_reg_psum_14_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_28( .activation_in(spare_reg_activation_14_27), .weight_in(spare_reg_weight_13_28), .partial_sum_in(spare_reg_psum_13_28), .reg_activation(spare_reg_activation_14_28), .reg_weight(spare_reg_weight_14_28), .reg_partial_sum(spare_reg_psum_14_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_29( .activation_in(spare_reg_activation_14_28), .weight_in(spare_reg_weight_13_29), .partial_sum_in(spare_reg_psum_13_29), .reg_activation(spare_reg_activation_14_29), .reg_weight(spare_reg_weight_14_29), .reg_partial_sum(spare_reg_psum_14_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_30( .activation_in(spare_reg_activation_14_29), .weight_in(spare_reg_weight_13_30), .partial_sum_in(spare_reg_psum_13_30), .reg_activation(spare_reg_activation_14_30), .reg_weight(spare_reg_weight_14_30), .reg_partial_sum(spare_reg_psum_14_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X14_31( .activation_in(spare_reg_activation_14_30), .weight_in(spare_reg_weight_13_31), .partial_sum_in(spare_reg_psum_13_31), .reg_weight(spare_reg_weight_14_31), .reg_partial_sum(spare_reg_psum_14_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_0( .activation_in(in_activation_15), .weight_in(spare_reg_weight_14_0), .partial_sum_in(spare_reg_psum_14_0), .reg_activation(spare_reg_activation_15_0), .reg_weight(spare_reg_weight_15_0), .reg_partial_sum(spare_reg_psum_15_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_1( .activation_in(spare_reg_activation_15_0), .weight_in(spare_reg_weight_14_1), .partial_sum_in(spare_reg_psum_14_1), .reg_activation(spare_reg_activation_15_1), .reg_weight(spare_reg_weight_15_1), .reg_partial_sum(spare_reg_psum_15_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_2( .activation_in(spare_reg_activation_15_1), .weight_in(spare_reg_weight_14_2), .partial_sum_in(spare_reg_psum_14_2), .reg_activation(spare_reg_activation_15_2), .reg_weight(spare_reg_weight_15_2), .reg_partial_sum(spare_reg_psum_15_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_3( .activation_in(spare_reg_activation_15_2), .weight_in(spare_reg_weight_14_3), .partial_sum_in(spare_reg_psum_14_3), .reg_activation(spare_reg_activation_15_3), .reg_weight(spare_reg_weight_15_3), .reg_partial_sum(spare_reg_psum_15_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_4( .activation_in(spare_reg_activation_15_3), .weight_in(spare_reg_weight_14_4), .partial_sum_in(spare_reg_psum_14_4), .reg_activation(spare_reg_activation_15_4), .reg_weight(spare_reg_weight_15_4), .reg_partial_sum(spare_reg_psum_15_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_5( .activation_in(spare_reg_activation_15_4), .weight_in(spare_reg_weight_14_5), .partial_sum_in(spare_reg_psum_14_5), .reg_activation(spare_reg_activation_15_5), .reg_weight(spare_reg_weight_15_5), .reg_partial_sum(spare_reg_psum_15_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_6( .activation_in(spare_reg_activation_15_5), .weight_in(spare_reg_weight_14_6), .partial_sum_in(spare_reg_psum_14_6), .reg_activation(spare_reg_activation_15_6), .reg_weight(spare_reg_weight_15_6), .reg_partial_sum(spare_reg_psum_15_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_7( .activation_in(spare_reg_activation_15_6), .weight_in(spare_reg_weight_14_7), .partial_sum_in(spare_reg_psum_14_7), .reg_activation(spare_reg_activation_15_7), .reg_weight(spare_reg_weight_15_7), .reg_partial_sum(spare_reg_psum_15_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_8( .activation_in(spare_reg_activation_15_7), .weight_in(spare_reg_weight_14_8), .partial_sum_in(spare_reg_psum_14_8), .reg_activation(spare_reg_activation_15_8), .reg_weight(spare_reg_weight_15_8), .reg_partial_sum(spare_reg_psum_15_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_9( .activation_in(spare_reg_activation_15_8), .weight_in(spare_reg_weight_14_9), .partial_sum_in(spare_reg_psum_14_9), .reg_activation(spare_reg_activation_15_9), .reg_weight(spare_reg_weight_15_9), .reg_partial_sum(spare_reg_psum_15_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_10( .activation_in(spare_reg_activation_15_9), .weight_in(spare_reg_weight_14_10), .partial_sum_in(spare_reg_psum_14_10), .reg_activation(spare_reg_activation_15_10), .reg_weight(spare_reg_weight_15_10), .reg_partial_sum(spare_reg_psum_15_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_11( .activation_in(spare_reg_activation_15_10), .weight_in(spare_reg_weight_14_11), .partial_sum_in(spare_reg_psum_14_11), .reg_activation(spare_reg_activation_15_11), .reg_weight(spare_reg_weight_15_11), .reg_partial_sum(spare_reg_psum_15_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_12( .activation_in(spare_reg_activation_15_11), .weight_in(spare_reg_weight_14_12), .partial_sum_in(spare_reg_psum_14_12), .reg_activation(spare_reg_activation_15_12), .reg_weight(spare_reg_weight_15_12), .reg_partial_sum(spare_reg_psum_15_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_13( .activation_in(spare_reg_activation_15_12), .weight_in(spare_reg_weight_14_13), .partial_sum_in(spare_reg_psum_14_13), .reg_activation(spare_reg_activation_15_13), .reg_weight(spare_reg_weight_15_13), .reg_partial_sum(spare_reg_psum_15_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_14( .activation_in(spare_reg_activation_15_13), .weight_in(spare_reg_weight_14_14), .partial_sum_in(spare_reg_psum_14_14), .reg_activation(spare_reg_activation_15_14), .reg_weight(spare_reg_weight_15_14), .reg_partial_sum(spare_reg_psum_15_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_15( .activation_in(spare_reg_activation_15_14), .weight_in(spare_reg_weight_14_15), .partial_sum_in(spare_reg_psum_14_15), .reg_activation(spare_reg_activation_15_15), .reg_weight(spare_reg_weight_15_15), .reg_partial_sum(spare_reg_psum_15_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_16( .activation_in(spare_reg_activation_15_15), .weight_in(spare_reg_weight_14_16), .partial_sum_in(spare_reg_psum_14_16), .reg_activation(spare_reg_activation_15_16), .reg_weight(spare_reg_weight_15_16), .reg_partial_sum(spare_reg_psum_15_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_17( .activation_in(spare_reg_activation_15_16), .weight_in(spare_reg_weight_14_17), .partial_sum_in(spare_reg_psum_14_17), .reg_activation(spare_reg_activation_15_17), .reg_weight(spare_reg_weight_15_17), .reg_partial_sum(spare_reg_psum_15_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_18( .activation_in(spare_reg_activation_15_17), .weight_in(spare_reg_weight_14_18), .partial_sum_in(spare_reg_psum_14_18), .reg_activation(spare_reg_activation_15_18), .reg_weight(spare_reg_weight_15_18), .reg_partial_sum(spare_reg_psum_15_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_19( .activation_in(spare_reg_activation_15_18), .weight_in(spare_reg_weight_14_19), .partial_sum_in(spare_reg_psum_14_19), .reg_activation(spare_reg_activation_15_19), .reg_weight(spare_reg_weight_15_19), .reg_partial_sum(spare_reg_psum_15_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_20( .activation_in(spare_reg_activation_15_19), .weight_in(spare_reg_weight_14_20), .partial_sum_in(spare_reg_psum_14_20), .reg_activation(spare_reg_activation_15_20), .reg_weight(spare_reg_weight_15_20), .reg_partial_sum(spare_reg_psum_15_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_21( .activation_in(spare_reg_activation_15_20), .weight_in(spare_reg_weight_14_21), .partial_sum_in(spare_reg_psum_14_21), .reg_activation(spare_reg_activation_15_21), .reg_weight(spare_reg_weight_15_21), .reg_partial_sum(spare_reg_psum_15_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_22( .activation_in(spare_reg_activation_15_21), .weight_in(spare_reg_weight_14_22), .partial_sum_in(spare_reg_psum_14_22), .reg_activation(spare_reg_activation_15_22), .reg_weight(spare_reg_weight_15_22), .reg_partial_sum(spare_reg_psum_15_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_23( .activation_in(spare_reg_activation_15_22), .weight_in(spare_reg_weight_14_23), .partial_sum_in(spare_reg_psum_14_23), .reg_activation(spare_reg_activation_15_23), .reg_weight(spare_reg_weight_15_23), .reg_partial_sum(spare_reg_psum_15_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_24( .activation_in(spare_reg_activation_15_23), .weight_in(spare_reg_weight_14_24), .partial_sum_in(spare_reg_psum_14_24), .reg_activation(spare_reg_activation_15_24), .reg_weight(spare_reg_weight_15_24), .reg_partial_sum(spare_reg_psum_15_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_25( .activation_in(spare_reg_activation_15_24), .weight_in(spare_reg_weight_14_25), .partial_sum_in(spare_reg_psum_14_25), .reg_activation(spare_reg_activation_15_25), .reg_weight(spare_reg_weight_15_25), .reg_partial_sum(spare_reg_psum_15_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_26( .activation_in(spare_reg_activation_15_25), .weight_in(spare_reg_weight_14_26), .partial_sum_in(spare_reg_psum_14_26), .reg_activation(spare_reg_activation_15_26), .reg_weight(spare_reg_weight_15_26), .reg_partial_sum(spare_reg_psum_15_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_27( .activation_in(spare_reg_activation_15_26), .weight_in(spare_reg_weight_14_27), .partial_sum_in(spare_reg_psum_14_27), .reg_activation(spare_reg_activation_15_27), .reg_weight(spare_reg_weight_15_27), .reg_partial_sum(spare_reg_psum_15_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_28( .activation_in(spare_reg_activation_15_27), .weight_in(spare_reg_weight_14_28), .partial_sum_in(spare_reg_psum_14_28), .reg_activation(spare_reg_activation_15_28), .reg_weight(spare_reg_weight_15_28), .reg_partial_sum(spare_reg_psum_15_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_29( .activation_in(spare_reg_activation_15_28), .weight_in(spare_reg_weight_14_29), .partial_sum_in(spare_reg_psum_14_29), .reg_activation(spare_reg_activation_15_29), .reg_weight(spare_reg_weight_15_29), .reg_partial_sum(spare_reg_psum_15_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_30( .activation_in(spare_reg_activation_15_29), .weight_in(spare_reg_weight_14_30), .partial_sum_in(spare_reg_psum_14_30), .reg_activation(spare_reg_activation_15_30), .reg_weight(spare_reg_weight_15_30), .reg_partial_sum(spare_reg_psum_15_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X15_31( .activation_in(spare_reg_activation_15_30), .weight_in(spare_reg_weight_14_31), .partial_sum_in(spare_reg_psum_14_31), .reg_weight(spare_reg_weight_15_31), .reg_partial_sum(spare_reg_psum_15_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_0( .activation_in(in_activation_16), .weight_in(spare_reg_weight_15_0), .partial_sum_in(spare_reg_psum_15_0), .reg_activation(spare_reg_activation_16_0), .reg_weight(spare_reg_weight_16_0), .reg_partial_sum(spare_reg_psum_16_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_1( .activation_in(spare_reg_activation_16_0), .weight_in(spare_reg_weight_15_1), .partial_sum_in(spare_reg_psum_15_1), .reg_activation(spare_reg_activation_16_1), .reg_weight(spare_reg_weight_16_1), .reg_partial_sum(spare_reg_psum_16_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_2( .activation_in(spare_reg_activation_16_1), .weight_in(spare_reg_weight_15_2), .partial_sum_in(spare_reg_psum_15_2), .reg_activation(spare_reg_activation_16_2), .reg_weight(spare_reg_weight_16_2), .reg_partial_sum(spare_reg_psum_16_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_3( .activation_in(spare_reg_activation_16_2), .weight_in(spare_reg_weight_15_3), .partial_sum_in(spare_reg_psum_15_3), .reg_activation(spare_reg_activation_16_3), .reg_weight(spare_reg_weight_16_3), .reg_partial_sum(spare_reg_psum_16_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_4( .activation_in(spare_reg_activation_16_3), .weight_in(spare_reg_weight_15_4), .partial_sum_in(spare_reg_psum_15_4), .reg_activation(spare_reg_activation_16_4), .reg_weight(spare_reg_weight_16_4), .reg_partial_sum(spare_reg_psum_16_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_5( .activation_in(spare_reg_activation_16_4), .weight_in(spare_reg_weight_15_5), .partial_sum_in(spare_reg_psum_15_5), .reg_activation(spare_reg_activation_16_5), .reg_weight(spare_reg_weight_16_5), .reg_partial_sum(spare_reg_psum_16_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_6( .activation_in(spare_reg_activation_16_5), .weight_in(spare_reg_weight_15_6), .partial_sum_in(spare_reg_psum_15_6), .reg_activation(spare_reg_activation_16_6), .reg_weight(spare_reg_weight_16_6), .reg_partial_sum(spare_reg_psum_16_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_7( .activation_in(spare_reg_activation_16_6), .weight_in(spare_reg_weight_15_7), .partial_sum_in(spare_reg_psum_15_7), .reg_activation(spare_reg_activation_16_7), .reg_weight(spare_reg_weight_16_7), .reg_partial_sum(spare_reg_psum_16_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_8( .activation_in(spare_reg_activation_16_7), .weight_in(spare_reg_weight_15_8), .partial_sum_in(spare_reg_psum_15_8), .reg_activation(spare_reg_activation_16_8), .reg_weight(spare_reg_weight_16_8), .reg_partial_sum(spare_reg_psum_16_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_9( .activation_in(spare_reg_activation_16_8), .weight_in(spare_reg_weight_15_9), .partial_sum_in(spare_reg_psum_15_9), .reg_activation(spare_reg_activation_16_9), .reg_weight(spare_reg_weight_16_9), .reg_partial_sum(spare_reg_psum_16_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_10( .activation_in(spare_reg_activation_16_9), .weight_in(spare_reg_weight_15_10), .partial_sum_in(spare_reg_psum_15_10), .reg_activation(spare_reg_activation_16_10), .reg_weight(spare_reg_weight_16_10), .reg_partial_sum(spare_reg_psum_16_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_11( .activation_in(spare_reg_activation_16_10), .weight_in(spare_reg_weight_15_11), .partial_sum_in(spare_reg_psum_15_11), .reg_activation(spare_reg_activation_16_11), .reg_weight(spare_reg_weight_16_11), .reg_partial_sum(spare_reg_psum_16_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_12( .activation_in(spare_reg_activation_16_11), .weight_in(spare_reg_weight_15_12), .partial_sum_in(spare_reg_psum_15_12), .reg_activation(spare_reg_activation_16_12), .reg_weight(spare_reg_weight_16_12), .reg_partial_sum(spare_reg_psum_16_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_13( .activation_in(spare_reg_activation_16_12), .weight_in(spare_reg_weight_15_13), .partial_sum_in(spare_reg_psum_15_13), .reg_activation(spare_reg_activation_16_13), .reg_weight(spare_reg_weight_16_13), .reg_partial_sum(spare_reg_psum_16_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_14( .activation_in(spare_reg_activation_16_13), .weight_in(spare_reg_weight_15_14), .partial_sum_in(spare_reg_psum_15_14), .reg_activation(spare_reg_activation_16_14), .reg_weight(spare_reg_weight_16_14), .reg_partial_sum(spare_reg_psum_16_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_15( .activation_in(spare_reg_activation_16_14), .weight_in(spare_reg_weight_15_15), .partial_sum_in(spare_reg_psum_15_15), .reg_activation(spare_reg_activation_16_15), .reg_weight(spare_reg_weight_16_15), .reg_partial_sum(spare_reg_psum_16_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_16( .activation_in(spare_reg_activation_16_15), .weight_in(spare_reg_weight_15_16), .partial_sum_in(spare_reg_psum_15_16), .reg_activation(spare_reg_activation_16_16), .reg_weight(spare_reg_weight_16_16), .reg_partial_sum(spare_reg_psum_16_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_17( .activation_in(spare_reg_activation_16_16), .weight_in(spare_reg_weight_15_17), .partial_sum_in(spare_reg_psum_15_17), .reg_activation(spare_reg_activation_16_17), .reg_weight(spare_reg_weight_16_17), .reg_partial_sum(spare_reg_psum_16_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_18( .activation_in(spare_reg_activation_16_17), .weight_in(spare_reg_weight_15_18), .partial_sum_in(spare_reg_psum_15_18), .reg_activation(spare_reg_activation_16_18), .reg_weight(spare_reg_weight_16_18), .reg_partial_sum(spare_reg_psum_16_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_19( .activation_in(spare_reg_activation_16_18), .weight_in(spare_reg_weight_15_19), .partial_sum_in(spare_reg_psum_15_19), .reg_activation(spare_reg_activation_16_19), .reg_weight(spare_reg_weight_16_19), .reg_partial_sum(spare_reg_psum_16_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_20( .activation_in(spare_reg_activation_16_19), .weight_in(spare_reg_weight_15_20), .partial_sum_in(spare_reg_psum_15_20), .reg_activation(spare_reg_activation_16_20), .reg_weight(spare_reg_weight_16_20), .reg_partial_sum(spare_reg_psum_16_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_21( .activation_in(spare_reg_activation_16_20), .weight_in(spare_reg_weight_15_21), .partial_sum_in(spare_reg_psum_15_21), .reg_activation(spare_reg_activation_16_21), .reg_weight(spare_reg_weight_16_21), .reg_partial_sum(spare_reg_psum_16_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_22( .activation_in(spare_reg_activation_16_21), .weight_in(spare_reg_weight_15_22), .partial_sum_in(spare_reg_psum_15_22), .reg_activation(spare_reg_activation_16_22), .reg_weight(spare_reg_weight_16_22), .reg_partial_sum(spare_reg_psum_16_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_23( .activation_in(spare_reg_activation_16_22), .weight_in(spare_reg_weight_15_23), .partial_sum_in(spare_reg_psum_15_23), .reg_activation(spare_reg_activation_16_23), .reg_weight(spare_reg_weight_16_23), .reg_partial_sum(spare_reg_psum_16_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_24( .activation_in(spare_reg_activation_16_23), .weight_in(spare_reg_weight_15_24), .partial_sum_in(spare_reg_psum_15_24), .reg_activation(spare_reg_activation_16_24), .reg_weight(spare_reg_weight_16_24), .reg_partial_sum(spare_reg_psum_16_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_25( .activation_in(spare_reg_activation_16_24), .weight_in(spare_reg_weight_15_25), .partial_sum_in(spare_reg_psum_15_25), .reg_activation(spare_reg_activation_16_25), .reg_weight(spare_reg_weight_16_25), .reg_partial_sum(spare_reg_psum_16_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_26( .activation_in(spare_reg_activation_16_25), .weight_in(spare_reg_weight_15_26), .partial_sum_in(spare_reg_psum_15_26), .reg_activation(spare_reg_activation_16_26), .reg_weight(spare_reg_weight_16_26), .reg_partial_sum(spare_reg_psum_16_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_27( .activation_in(spare_reg_activation_16_26), .weight_in(spare_reg_weight_15_27), .partial_sum_in(spare_reg_psum_15_27), .reg_activation(spare_reg_activation_16_27), .reg_weight(spare_reg_weight_16_27), .reg_partial_sum(spare_reg_psum_16_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_28( .activation_in(spare_reg_activation_16_27), .weight_in(spare_reg_weight_15_28), .partial_sum_in(spare_reg_psum_15_28), .reg_activation(spare_reg_activation_16_28), .reg_weight(spare_reg_weight_16_28), .reg_partial_sum(spare_reg_psum_16_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_29( .activation_in(spare_reg_activation_16_28), .weight_in(spare_reg_weight_15_29), .partial_sum_in(spare_reg_psum_15_29), .reg_activation(spare_reg_activation_16_29), .reg_weight(spare_reg_weight_16_29), .reg_partial_sum(spare_reg_psum_16_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_30( .activation_in(spare_reg_activation_16_29), .weight_in(spare_reg_weight_15_30), .partial_sum_in(spare_reg_psum_15_30), .reg_activation(spare_reg_activation_16_30), .reg_weight(spare_reg_weight_16_30), .reg_partial_sum(spare_reg_psum_16_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X16_31( .activation_in(spare_reg_activation_16_30), .weight_in(spare_reg_weight_15_31), .partial_sum_in(spare_reg_psum_15_31), .reg_weight(spare_reg_weight_16_31), .reg_partial_sum(spare_reg_psum_16_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_0( .activation_in(in_activation_17), .weight_in(spare_reg_weight_16_0), .partial_sum_in(spare_reg_psum_16_0), .reg_activation(spare_reg_activation_17_0), .reg_weight(spare_reg_weight_17_0), .reg_partial_sum(spare_reg_psum_17_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_1( .activation_in(spare_reg_activation_17_0), .weight_in(spare_reg_weight_16_1), .partial_sum_in(spare_reg_psum_16_1), .reg_activation(spare_reg_activation_17_1), .reg_weight(spare_reg_weight_17_1), .reg_partial_sum(spare_reg_psum_17_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_2( .activation_in(spare_reg_activation_17_1), .weight_in(spare_reg_weight_16_2), .partial_sum_in(spare_reg_psum_16_2), .reg_activation(spare_reg_activation_17_2), .reg_weight(spare_reg_weight_17_2), .reg_partial_sum(spare_reg_psum_17_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_3( .activation_in(spare_reg_activation_17_2), .weight_in(spare_reg_weight_16_3), .partial_sum_in(spare_reg_psum_16_3), .reg_activation(spare_reg_activation_17_3), .reg_weight(spare_reg_weight_17_3), .reg_partial_sum(spare_reg_psum_17_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_4( .activation_in(spare_reg_activation_17_3), .weight_in(spare_reg_weight_16_4), .partial_sum_in(spare_reg_psum_16_4), .reg_activation(spare_reg_activation_17_4), .reg_weight(spare_reg_weight_17_4), .reg_partial_sum(spare_reg_psum_17_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_5( .activation_in(spare_reg_activation_17_4), .weight_in(spare_reg_weight_16_5), .partial_sum_in(spare_reg_psum_16_5), .reg_activation(spare_reg_activation_17_5), .reg_weight(spare_reg_weight_17_5), .reg_partial_sum(spare_reg_psum_17_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_6( .activation_in(spare_reg_activation_17_5), .weight_in(spare_reg_weight_16_6), .partial_sum_in(spare_reg_psum_16_6), .reg_activation(spare_reg_activation_17_6), .reg_weight(spare_reg_weight_17_6), .reg_partial_sum(spare_reg_psum_17_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_7( .activation_in(spare_reg_activation_17_6), .weight_in(spare_reg_weight_16_7), .partial_sum_in(spare_reg_psum_16_7), .reg_activation(spare_reg_activation_17_7), .reg_weight(spare_reg_weight_17_7), .reg_partial_sum(spare_reg_psum_17_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_8( .activation_in(spare_reg_activation_17_7), .weight_in(spare_reg_weight_16_8), .partial_sum_in(spare_reg_psum_16_8), .reg_activation(spare_reg_activation_17_8), .reg_weight(spare_reg_weight_17_8), .reg_partial_sum(spare_reg_psum_17_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_9( .activation_in(spare_reg_activation_17_8), .weight_in(spare_reg_weight_16_9), .partial_sum_in(spare_reg_psum_16_9), .reg_activation(spare_reg_activation_17_9), .reg_weight(spare_reg_weight_17_9), .reg_partial_sum(spare_reg_psum_17_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_10( .activation_in(spare_reg_activation_17_9), .weight_in(spare_reg_weight_16_10), .partial_sum_in(spare_reg_psum_16_10), .reg_activation(spare_reg_activation_17_10), .reg_weight(spare_reg_weight_17_10), .reg_partial_sum(spare_reg_psum_17_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_11( .activation_in(spare_reg_activation_17_10), .weight_in(spare_reg_weight_16_11), .partial_sum_in(spare_reg_psum_16_11), .reg_activation(spare_reg_activation_17_11), .reg_weight(spare_reg_weight_17_11), .reg_partial_sum(spare_reg_psum_17_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_12( .activation_in(spare_reg_activation_17_11), .weight_in(spare_reg_weight_16_12), .partial_sum_in(spare_reg_psum_16_12), .reg_activation(spare_reg_activation_17_12), .reg_weight(spare_reg_weight_17_12), .reg_partial_sum(spare_reg_psum_17_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_13( .activation_in(spare_reg_activation_17_12), .weight_in(spare_reg_weight_16_13), .partial_sum_in(spare_reg_psum_16_13), .reg_activation(spare_reg_activation_17_13), .reg_weight(spare_reg_weight_17_13), .reg_partial_sum(spare_reg_psum_17_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_14( .activation_in(spare_reg_activation_17_13), .weight_in(spare_reg_weight_16_14), .partial_sum_in(spare_reg_psum_16_14), .reg_activation(spare_reg_activation_17_14), .reg_weight(spare_reg_weight_17_14), .reg_partial_sum(spare_reg_psum_17_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_15( .activation_in(spare_reg_activation_17_14), .weight_in(spare_reg_weight_16_15), .partial_sum_in(spare_reg_psum_16_15), .reg_activation(spare_reg_activation_17_15), .reg_weight(spare_reg_weight_17_15), .reg_partial_sum(spare_reg_psum_17_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_16( .activation_in(spare_reg_activation_17_15), .weight_in(spare_reg_weight_16_16), .partial_sum_in(spare_reg_psum_16_16), .reg_activation(spare_reg_activation_17_16), .reg_weight(spare_reg_weight_17_16), .reg_partial_sum(spare_reg_psum_17_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_17( .activation_in(spare_reg_activation_17_16), .weight_in(spare_reg_weight_16_17), .partial_sum_in(spare_reg_psum_16_17), .reg_activation(spare_reg_activation_17_17), .reg_weight(spare_reg_weight_17_17), .reg_partial_sum(spare_reg_psum_17_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_18( .activation_in(spare_reg_activation_17_17), .weight_in(spare_reg_weight_16_18), .partial_sum_in(spare_reg_psum_16_18), .reg_activation(spare_reg_activation_17_18), .reg_weight(spare_reg_weight_17_18), .reg_partial_sum(spare_reg_psum_17_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_19( .activation_in(spare_reg_activation_17_18), .weight_in(spare_reg_weight_16_19), .partial_sum_in(spare_reg_psum_16_19), .reg_activation(spare_reg_activation_17_19), .reg_weight(spare_reg_weight_17_19), .reg_partial_sum(spare_reg_psum_17_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_20( .activation_in(spare_reg_activation_17_19), .weight_in(spare_reg_weight_16_20), .partial_sum_in(spare_reg_psum_16_20), .reg_activation(spare_reg_activation_17_20), .reg_weight(spare_reg_weight_17_20), .reg_partial_sum(spare_reg_psum_17_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_21( .activation_in(spare_reg_activation_17_20), .weight_in(spare_reg_weight_16_21), .partial_sum_in(spare_reg_psum_16_21), .reg_activation(spare_reg_activation_17_21), .reg_weight(spare_reg_weight_17_21), .reg_partial_sum(spare_reg_psum_17_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_22( .activation_in(spare_reg_activation_17_21), .weight_in(spare_reg_weight_16_22), .partial_sum_in(spare_reg_psum_16_22), .reg_activation(spare_reg_activation_17_22), .reg_weight(spare_reg_weight_17_22), .reg_partial_sum(spare_reg_psum_17_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_23( .activation_in(spare_reg_activation_17_22), .weight_in(spare_reg_weight_16_23), .partial_sum_in(spare_reg_psum_16_23), .reg_activation(spare_reg_activation_17_23), .reg_weight(spare_reg_weight_17_23), .reg_partial_sum(spare_reg_psum_17_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_24( .activation_in(spare_reg_activation_17_23), .weight_in(spare_reg_weight_16_24), .partial_sum_in(spare_reg_psum_16_24), .reg_activation(spare_reg_activation_17_24), .reg_weight(spare_reg_weight_17_24), .reg_partial_sum(spare_reg_psum_17_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_25( .activation_in(spare_reg_activation_17_24), .weight_in(spare_reg_weight_16_25), .partial_sum_in(spare_reg_psum_16_25), .reg_activation(spare_reg_activation_17_25), .reg_weight(spare_reg_weight_17_25), .reg_partial_sum(spare_reg_psum_17_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_26( .activation_in(spare_reg_activation_17_25), .weight_in(spare_reg_weight_16_26), .partial_sum_in(spare_reg_psum_16_26), .reg_activation(spare_reg_activation_17_26), .reg_weight(spare_reg_weight_17_26), .reg_partial_sum(spare_reg_psum_17_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_27( .activation_in(spare_reg_activation_17_26), .weight_in(spare_reg_weight_16_27), .partial_sum_in(spare_reg_psum_16_27), .reg_activation(spare_reg_activation_17_27), .reg_weight(spare_reg_weight_17_27), .reg_partial_sum(spare_reg_psum_17_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_28( .activation_in(spare_reg_activation_17_27), .weight_in(spare_reg_weight_16_28), .partial_sum_in(spare_reg_psum_16_28), .reg_activation(spare_reg_activation_17_28), .reg_weight(spare_reg_weight_17_28), .reg_partial_sum(spare_reg_psum_17_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_29( .activation_in(spare_reg_activation_17_28), .weight_in(spare_reg_weight_16_29), .partial_sum_in(spare_reg_psum_16_29), .reg_activation(spare_reg_activation_17_29), .reg_weight(spare_reg_weight_17_29), .reg_partial_sum(spare_reg_psum_17_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_30( .activation_in(spare_reg_activation_17_29), .weight_in(spare_reg_weight_16_30), .partial_sum_in(spare_reg_psum_16_30), .reg_activation(spare_reg_activation_17_30), .reg_weight(spare_reg_weight_17_30), .reg_partial_sum(spare_reg_psum_17_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X17_31( .activation_in(spare_reg_activation_17_30), .weight_in(spare_reg_weight_16_31), .partial_sum_in(spare_reg_psum_16_31), .reg_weight(spare_reg_weight_17_31), .reg_partial_sum(spare_reg_psum_17_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_0( .activation_in(in_activation_18), .weight_in(spare_reg_weight_17_0), .partial_sum_in(spare_reg_psum_17_0), .reg_activation(spare_reg_activation_18_0), .reg_weight(spare_reg_weight_18_0), .reg_partial_sum(spare_reg_psum_18_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_1( .activation_in(spare_reg_activation_18_0), .weight_in(spare_reg_weight_17_1), .partial_sum_in(spare_reg_psum_17_1), .reg_activation(spare_reg_activation_18_1), .reg_weight(spare_reg_weight_18_1), .reg_partial_sum(spare_reg_psum_18_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_2( .activation_in(spare_reg_activation_18_1), .weight_in(spare_reg_weight_17_2), .partial_sum_in(spare_reg_psum_17_2), .reg_activation(spare_reg_activation_18_2), .reg_weight(spare_reg_weight_18_2), .reg_partial_sum(spare_reg_psum_18_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_3( .activation_in(spare_reg_activation_18_2), .weight_in(spare_reg_weight_17_3), .partial_sum_in(spare_reg_psum_17_3), .reg_activation(spare_reg_activation_18_3), .reg_weight(spare_reg_weight_18_3), .reg_partial_sum(spare_reg_psum_18_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_4( .activation_in(spare_reg_activation_18_3), .weight_in(spare_reg_weight_17_4), .partial_sum_in(spare_reg_psum_17_4), .reg_activation(spare_reg_activation_18_4), .reg_weight(spare_reg_weight_18_4), .reg_partial_sum(spare_reg_psum_18_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_5( .activation_in(spare_reg_activation_18_4), .weight_in(spare_reg_weight_17_5), .partial_sum_in(spare_reg_psum_17_5), .reg_activation(spare_reg_activation_18_5), .reg_weight(spare_reg_weight_18_5), .reg_partial_sum(spare_reg_psum_18_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_6( .activation_in(spare_reg_activation_18_5), .weight_in(spare_reg_weight_17_6), .partial_sum_in(spare_reg_psum_17_6), .reg_activation(spare_reg_activation_18_6), .reg_weight(spare_reg_weight_18_6), .reg_partial_sum(spare_reg_psum_18_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_7( .activation_in(spare_reg_activation_18_6), .weight_in(spare_reg_weight_17_7), .partial_sum_in(spare_reg_psum_17_7), .reg_activation(spare_reg_activation_18_7), .reg_weight(spare_reg_weight_18_7), .reg_partial_sum(spare_reg_psum_18_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_8( .activation_in(spare_reg_activation_18_7), .weight_in(spare_reg_weight_17_8), .partial_sum_in(spare_reg_psum_17_8), .reg_activation(spare_reg_activation_18_8), .reg_weight(spare_reg_weight_18_8), .reg_partial_sum(spare_reg_psum_18_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_9( .activation_in(spare_reg_activation_18_8), .weight_in(spare_reg_weight_17_9), .partial_sum_in(spare_reg_psum_17_9), .reg_activation(spare_reg_activation_18_9), .reg_weight(spare_reg_weight_18_9), .reg_partial_sum(spare_reg_psum_18_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_10( .activation_in(spare_reg_activation_18_9), .weight_in(spare_reg_weight_17_10), .partial_sum_in(spare_reg_psum_17_10), .reg_activation(spare_reg_activation_18_10), .reg_weight(spare_reg_weight_18_10), .reg_partial_sum(spare_reg_psum_18_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_11( .activation_in(spare_reg_activation_18_10), .weight_in(spare_reg_weight_17_11), .partial_sum_in(spare_reg_psum_17_11), .reg_activation(spare_reg_activation_18_11), .reg_weight(spare_reg_weight_18_11), .reg_partial_sum(spare_reg_psum_18_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_12( .activation_in(spare_reg_activation_18_11), .weight_in(spare_reg_weight_17_12), .partial_sum_in(spare_reg_psum_17_12), .reg_activation(spare_reg_activation_18_12), .reg_weight(spare_reg_weight_18_12), .reg_partial_sum(spare_reg_psum_18_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_13( .activation_in(spare_reg_activation_18_12), .weight_in(spare_reg_weight_17_13), .partial_sum_in(spare_reg_psum_17_13), .reg_activation(spare_reg_activation_18_13), .reg_weight(spare_reg_weight_18_13), .reg_partial_sum(spare_reg_psum_18_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_14( .activation_in(spare_reg_activation_18_13), .weight_in(spare_reg_weight_17_14), .partial_sum_in(spare_reg_psum_17_14), .reg_activation(spare_reg_activation_18_14), .reg_weight(spare_reg_weight_18_14), .reg_partial_sum(spare_reg_psum_18_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_15( .activation_in(spare_reg_activation_18_14), .weight_in(spare_reg_weight_17_15), .partial_sum_in(spare_reg_psum_17_15), .reg_activation(spare_reg_activation_18_15), .reg_weight(spare_reg_weight_18_15), .reg_partial_sum(spare_reg_psum_18_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_16( .activation_in(spare_reg_activation_18_15), .weight_in(spare_reg_weight_17_16), .partial_sum_in(spare_reg_psum_17_16), .reg_activation(spare_reg_activation_18_16), .reg_weight(spare_reg_weight_18_16), .reg_partial_sum(spare_reg_psum_18_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_17( .activation_in(spare_reg_activation_18_16), .weight_in(spare_reg_weight_17_17), .partial_sum_in(spare_reg_psum_17_17), .reg_activation(spare_reg_activation_18_17), .reg_weight(spare_reg_weight_18_17), .reg_partial_sum(spare_reg_psum_18_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_18( .activation_in(spare_reg_activation_18_17), .weight_in(spare_reg_weight_17_18), .partial_sum_in(spare_reg_psum_17_18), .reg_activation(spare_reg_activation_18_18), .reg_weight(spare_reg_weight_18_18), .reg_partial_sum(spare_reg_psum_18_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_19( .activation_in(spare_reg_activation_18_18), .weight_in(spare_reg_weight_17_19), .partial_sum_in(spare_reg_psum_17_19), .reg_activation(spare_reg_activation_18_19), .reg_weight(spare_reg_weight_18_19), .reg_partial_sum(spare_reg_psum_18_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_20( .activation_in(spare_reg_activation_18_19), .weight_in(spare_reg_weight_17_20), .partial_sum_in(spare_reg_psum_17_20), .reg_activation(spare_reg_activation_18_20), .reg_weight(spare_reg_weight_18_20), .reg_partial_sum(spare_reg_psum_18_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_21( .activation_in(spare_reg_activation_18_20), .weight_in(spare_reg_weight_17_21), .partial_sum_in(spare_reg_psum_17_21), .reg_activation(spare_reg_activation_18_21), .reg_weight(spare_reg_weight_18_21), .reg_partial_sum(spare_reg_psum_18_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_22( .activation_in(spare_reg_activation_18_21), .weight_in(spare_reg_weight_17_22), .partial_sum_in(spare_reg_psum_17_22), .reg_activation(spare_reg_activation_18_22), .reg_weight(spare_reg_weight_18_22), .reg_partial_sum(spare_reg_psum_18_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_23( .activation_in(spare_reg_activation_18_22), .weight_in(spare_reg_weight_17_23), .partial_sum_in(spare_reg_psum_17_23), .reg_activation(spare_reg_activation_18_23), .reg_weight(spare_reg_weight_18_23), .reg_partial_sum(spare_reg_psum_18_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_24( .activation_in(spare_reg_activation_18_23), .weight_in(spare_reg_weight_17_24), .partial_sum_in(spare_reg_psum_17_24), .reg_activation(spare_reg_activation_18_24), .reg_weight(spare_reg_weight_18_24), .reg_partial_sum(spare_reg_psum_18_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_25( .activation_in(spare_reg_activation_18_24), .weight_in(spare_reg_weight_17_25), .partial_sum_in(spare_reg_psum_17_25), .reg_activation(spare_reg_activation_18_25), .reg_weight(spare_reg_weight_18_25), .reg_partial_sum(spare_reg_psum_18_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_26( .activation_in(spare_reg_activation_18_25), .weight_in(spare_reg_weight_17_26), .partial_sum_in(spare_reg_psum_17_26), .reg_activation(spare_reg_activation_18_26), .reg_weight(spare_reg_weight_18_26), .reg_partial_sum(spare_reg_psum_18_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_27( .activation_in(spare_reg_activation_18_26), .weight_in(spare_reg_weight_17_27), .partial_sum_in(spare_reg_psum_17_27), .reg_activation(spare_reg_activation_18_27), .reg_weight(spare_reg_weight_18_27), .reg_partial_sum(spare_reg_psum_18_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_28( .activation_in(spare_reg_activation_18_27), .weight_in(spare_reg_weight_17_28), .partial_sum_in(spare_reg_psum_17_28), .reg_activation(spare_reg_activation_18_28), .reg_weight(spare_reg_weight_18_28), .reg_partial_sum(spare_reg_psum_18_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_29( .activation_in(spare_reg_activation_18_28), .weight_in(spare_reg_weight_17_29), .partial_sum_in(spare_reg_psum_17_29), .reg_activation(spare_reg_activation_18_29), .reg_weight(spare_reg_weight_18_29), .reg_partial_sum(spare_reg_psum_18_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_30( .activation_in(spare_reg_activation_18_29), .weight_in(spare_reg_weight_17_30), .partial_sum_in(spare_reg_psum_17_30), .reg_activation(spare_reg_activation_18_30), .reg_weight(spare_reg_weight_18_30), .reg_partial_sum(spare_reg_psum_18_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X18_31( .activation_in(spare_reg_activation_18_30), .weight_in(spare_reg_weight_17_31), .partial_sum_in(spare_reg_psum_17_31), .reg_weight(spare_reg_weight_18_31), .reg_partial_sum(spare_reg_psum_18_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_0( .activation_in(in_activation_19), .weight_in(spare_reg_weight_18_0), .partial_sum_in(spare_reg_psum_18_0), .reg_activation(spare_reg_activation_19_0), .reg_weight(spare_reg_weight_19_0), .reg_partial_sum(spare_reg_psum_19_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_1( .activation_in(spare_reg_activation_19_0), .weight_in(spare_reg_weight_18_1), .partial_sum_in(spare_reg_psum_18_1), .reg_activation(spare_reg_activation_19_1), .reg_weight(spare_reg_weight_19_1), .reg_partial_sum(spare_reg_psum_19_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_2( .activation_in(spare_reg_activation_19_1), .weight_in(spare_reg_weight_18_2), .partial_sum_in(spare_reg_psum_18_2), .reg_activation(spare_reg_activation_19_2), .reg_weight(spare_reg_weight_19_2), .reg_partial_sum(spare_reg_psum_19_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_3( .activation_in(spare_reg_activation_19_2), .weight_in(spare_reg_weight_18_3), .partial_sum_in(spare_reg_psum_18_3), .reg_activation(spare_reg_activation_19_3), .reg_weight(spare_reg_weight_19_3), .reg_partial_sum(spare_reg_psum_19_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_4( .activation_in(spare_reg_activation_19_3), .weight_in(spare_reg_weight_18_4), .partial_sum_in(spare_reg_psum_18_4), .reg_activation(spare_reg_activation_19_4), .reg_weight(spare_reg_weight_19_4), .reg_partial_sum(spare_reg_psum_19_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_5( .activation_in(spare_reg_activation_19_4), .weight_in(spare_reg_weight_18_5), .partial_sum_in(spare_reg_psum_18_5), .reg_activation(spare_reg_activation_19_5), .reg_weight(spare_reg_weight_19_5), .reg_partial_sum(spare_reg_psum_19_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_6( .activation_in(spare_reg_activation_19_5), .weight_in(spare_reg_weight_18_6), .partial_sum_in(spare_reg_psum_18_6), .reg_activation(spare_reg_activation_19_6), .reg_weight(spare_reg_weight_19_6), .reg_partial_sum(spare_reg_psum_19_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_7( .activation_in(spare_reg_activation_19_6), .weight_in(spare_reg_weight_18_7), .partial_sum_in(spare_reg_psum_18_7), .reg_activation(spare_reg_activation_19_7), .reg_weight(spare_reg_weight_19_7), .reg_partial_sum(spare_reg_psum_19_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_8( .activation_in(spare_reg_activation_19_7), .weight_in(spare_reg_weight_18_8), .partial_sum_in(spare_reg_psum_18_8), .reg_activation(spare_reg_activation_19_8), .reg_weight(spare_reg_weight_19_8), .reg_partial_sum(spare_reg_psum_19_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_9( .activation_in(spare_reg_activation_19_8), .weight_in(spare_reg_weight_18_9), .partial_sum_in(spare_reg_psum_18_9), .reg_activation(spare_reg_activation_19_9), .reg_weight(spare_reg_weight_19_9), .reg_partial_sum(spare_reg_psum_19_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_10( .activation_in(spare_reg_activation_19_9), .weight_in(spare_reg_weight_18_10), .partial_sum_in(spare_reg_psum_18_10), .reg_activation(spare_reg_activation_19_10), .reg_weight(spare_reg_weight_19_10), .reg_partial_sum(spare_reg_psum_19_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_11( .activation_in(spare_reg_activation_19_10), .weight_in(spare_reg_weight_18_11), .partial_sum_in(spare_reg_psum_18_11), .reg_activation(spare_reg_activation_19_11), .reg_weight(spare_reg_weight_19_11), .reg_partial_sum(spare_reg_psum_19_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_12( .activation_in(spare_reg_activation_19_11), .weight_in(spare_reg_weight_18_12), .partial_sum_in(spare_reg_psum_18_12), .reg_activation(spare_reg_activation_19_12), .reg_weight(spare_reg_weight_19_12), .reg_partial_sum(spare_reg_psum_19_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_13( .activation_in(spare_reg_activation_19_12), .weight_in(spare_reg_weight_18_13), .partial_sum_in(spare_reg_psum_18_13), .reg_activation(spare_reg_activation_19_13), .reg_weight(spare_reg_weight_19_13), .reg_partial_sum(spare_reg_psum_19_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_14( .activation_in(spare_reg_activation_19_13), .weight_in(spare_reg_weight_18_14), .partial_sum_in(spare_reg_psum_18_14), .reg_activation(spare_reg_activation_19_14), .reg_weight(spare_reg_weight_19_14), .reg_partial_sum(spare_reg_psum_19_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_15( .activation_in(spare_reg_activation_19_14), .weight_in(spare_reg_weight_18_15), .partial_sum_in(spare_reg_psum_18_15), .reg_activation(spare_reg_activation_19_15), .reg_weight(spare_reg_weight_19_15), .reg_partial_sum(spare_reg_psum_19_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_16( .activation_in(spare_reg_activation_19_15), .weight_in(spare_reg_weight_18_16), .partial_sum_in(spare_reg_psum_18_16), .reg_activation(spare_reg_activation_19_16), .reg_weight(spare_reg_weight_19_16), .reg_partial_sum(spare_reg_psum_19_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_17( .activation_in(spare_reg_activation_19_16), .weight_in(spare_reg_weight_18_17), .partial_sum_in(spare_reg_psum_18_17), .reg_activation(spare_reg_activation_19_17), .reg_weight(spare_reg_weight_19_17), .reg_partial_sum(spare_reg_psum_19_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_18( .activation_in(spare_reg_activation_19_17), .weight_in(spare_reg_weight_18_18), .partial_sum_in(spare_reg_psum_18_18), .reg_activation(spare_reg_activation_19_18), .reg_weight(spare_reg_weight_19_18), .reg_partial_sum(spare_reg_psum_19_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_19( .activation_in(spare_reg_activation_19_18), .weight_in(spare_reg_weight_18_19), .partial_sum_in(spare_reg_psum_18_19), .reg_activation(spare_reg_activation_19_19), .reg_weight(spare_reg_weight_19_19), .reg_partial_sum(spare_reg_psum_19_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_20( .activation_in(spare_reg_activation_19_19), .weight_in(spare_reg_weight_18_20), .partial_sum_in(spare_reg_psum_18_20), .reg_activation(spare_reg_activation_19_20), .reg_weight(spare_reg_weight_19_20), .reg_partial_sum(spare_reg_psum_19_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_21( .activation_in(spare_reg_activation_19_20), .weight_in(spare_reg_weight_18_21), .partial_sum_in(spare_reg_psum_18_21), .reg_activation(spare_reg_activation_19_21), .reg_weight(spare_reg_weight_19_21), .reg_partial_sum(spare_reg_psum_19_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_22( .activation_in(spare_reg_activation_19_21), .weight_in(spare_reg_weight_18_22), .partial_sum_in(spare_reg_psum_18_22), .reg_activation(spare_reg_activation_19_22), .reg_weight(spare_reg_weight_19_22), .reg_partial_sum(spare_reg_psum_19_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_23( .activation_in(spare_reg_activation_19_22), .weight_in(spare_reg_weight_18_23), .partial_sum_in(spare_reg_psum_18_23), .reg_activation(spare_reg_activation_19_23), .reg_weight(spare_reg_weight_19_23), .reg_partial_sum(spare_reg_psum_19_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_24( .activation_in(spare_reg_activation_19_23), .weight_in(spare_reg_weight_18_24), .partial_sum_in(spare_reg_psum_18_24), .reg_activation(spare_reg_activation_19_24), .reg_weight(spare_reg_weight_19_24), .reg_partial_sum(spare_reg_psum_19_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_25( .activation_in(spare_reg_activation_19_24), .weight_in(spare_reg_weight_18_25), .partial_sum_in(spare_reg_psum_18_25), .reg_activation(spare_reg_activation_19_25), .reg_weight(spare_reg_weight_19_25), .reg_partial_sum(spare_reg_psum_19_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_26( .activation_in(spare_reg_activation_19_25), .weight_in(spare_reg_weight_18_26), .partial_sum_in(spare_reg_psum_18_26), .reg_activation(spare_reg_activation_19_26), .reg_weight(spare_reg_weight_19_26), .reg_partial_sum(spare_reg_psum_19_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_27( .activation_in(spare_reg_activation_19_26), .weight_in(spare_reg_weight_18_27), .partial_sum_in(spare_reg_psum_18_27), .reg_activation(spare_reg_activation_19_27), .reg_weight(spare_reg_weight_19_27), .reg_partial_sum(spare_reg_psum_19_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_28( .activation_in(spare_reg_activation_19_27), .weight_in(spare_reg_weight_18_28), .partial_sum_in(spare_reg_psum_18_28), .reg_activation(spare_reg_activation_19_28), .reg_weight(spare_reg_weight_19_28), .reg_partial_sum(spare_reg_psum_19_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_29( .activation_in(spare_reg_activation_19_28), .weight_in(spare_reg_weight_18_29), .partial_sum_in(spare_reg_psum_18_29), .reg_activation(spare_reg_activation_19_29), .reg_weight(spare_reg_weight_19_29), .reg_partial_sum(spare_reg_psum_19_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_30( .activation_in(spare_reg_activation_19_29), .weight_in(spare_reg_weight_18_30), .partial_sum_in(spare_reg_psum_18_30), .reg_activation(spare_reg_activation_19_30), .reg_weight(spare_reg_weight_19_30), .reg_partial_sum(spare_reg_psum_19_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X19_31( .activation_in(spare_reg_activation_19_30), .weight_in(spare_reg_weight_18_31), .partial_sum_in(spare_reg_psum_18_31), .reg_weight(spare_reg_weight_19_31), .reg_partial_sum(spare_reg_psum_19_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_0( .activation_in(in_activation_20), .weight_in(spare_reg_weight_19_0), .partial_sum_in(spare_reg_psum_19_0), .reg_activation(spare_reg_activation_20_0), .reg_weight(spare_reg_weight_20_0), .reg_partial_sum(spare_reg_psum_20_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_1( .activation_in(spare_reg_activation_20_0), .weight_in(spare_reg_weight_19_1), .partial_sum_in(spare_reg_psum_19_1), .reg_activation(spare_reg_activation_20_1), .reg_weight(spare_reg_weight_20_1), .reg_partial_sum(spare_reg_psum_20_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_2( .activation_in(spare_reg_activation_20_1), .weight_in(spare_reg_weight_19_2), .partial_sum_in(spare_reg_psum_19_2), .reg_activation(spare_reg_activation_20_2), .reg_weight(spare_reg_weight_20_2), .reg_partial_sum(spare_reg_psum_20_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_3( .activation_in(spare_reg_activation_20_2), .weight_in(spare_reg_weight_19_3), .partial_sum_in(spare_reg_psum_19_3), .reg_activation(spare_reg_activation_20_3), .reg_weight(spare_reg_weight_20_3), .reg_partial_sum(spare_reg_psum_20_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_4( .activation_in(spare_reg_activation_20_3), .weight_in(spare_reg_weight_19_4), .partial_sum_in(spare_reg_psum_19_4), .reg_activation(spare_reg_activation_20_4), .reg_weight(spare_reg_weight_20_4), .reg_partial_sum(spare_reg_psum_20_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_5( .activation_in(spare_reg_activation_20_4), .weight_in(spare_reg_weight_19_5), .partial_sum_in(spare_reg_psum_19_5), .reg_activation(spare_reg_activation_20_5), .reg_weight(spare_reg_weight_20_5), .reg_partial_sum(spare_reg_psum_20_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_6( .activation_in(spare_reg_activation_20_5), .weight_in(spare_reg_weight_19_6), .partial_sum_in(spare_reg_psum_19_6), .reg_activation(spare_reg_activation_20_6), .reg_weight(spare_reg_weight_20_6), .reg_partial_sum(spare_reg_psum_20_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_7( .activation_in(spare_reg_activation_20_6), .weight_in(spare_reg_weight_19_7), .partial_sum_in(spare_reg_psum_19_7), .reg_activation(spare_reg_activation_20_7), .reg_weight(spare_reg_weight_20_7), .reg_partial_sum(spare_reg_psum_20_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_8( .activation_in(spare_reg_activation_20_7), .weight_in(spare_reg_weight_19_8), .partial_sum_in(spare_reg_psum_19_8), .reg_activation(spare_reg_activation_20_8), .reg_weight(spare_reg_weight_20_8), .reg_partial_sum(spare_reg_psum_20_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_9( .activation_in(spare_reg_activation_20_8), .weight_in(spare_reg_weight_19_9), .partial_sum_in(spare_reg_psum_19_9), .reg_activation(spare_reg_activation_20_9), .reg_weight(spare_reg_weight_20_9), .reg_partial_sum(spare_reg_psum_20_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_10( .activation_in(spare_reg_activation_20_9), .weight_in(spare_reg_weight_19_10), .partial_sum_in(spare_reg_psum_19_10), .reg_activation(spare_reg_activation_20_10), .reg_weight(spare_reg_weight_20_10), .reg_partial_sum(spare_reg_psum_20_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_11( .activation_in(spare_reg_activation_20_10), .weight_in(spare_reg_weight_19_11), .partial_sum_in(spare_reg_psum_19_11), .reg_activation(spare_reg_activation_20_11), .reg_weight(spare_reg_weight_20_11), .reg_partial_sum(spare_reg_psum_20_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_12( .activation_in(spare_reg_activation_20_11), .weight_in(spare_reg_weight_19_12), .partial_sum_in(spare_reg_psum_19_12), .reg_activation(spare_reg_activation_20_12), .reg_weight(spare_reg_weight_20_12), .reg_partial_sum(spare_reg_psum_20_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_13( .activation_in(spare_reg_activation_20_12), .weight_in(spare_reg_weight_19_13), .partial_sum_in(spare_reg_psum_19_13), .reg_activation(spare_reg_activation_20_13), .reg_weight(spare_reg_weight_20_13), .reg_partial_sum(spare_reg_psum_20_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_14( .activation_in(spare_reg_activation_20_13), .weight_in(spare_reg_weight_19_14), .partial_sum_in(spare_reg_psum_19_14), .reg_activation(spare_reg_activation_20_14), .reg_weight(spare_reg_weight_20_14), .reg_partial_sum(spare_reg_psum_20_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_15( .activation_in(spare_reg_activation_20_14), .weight_in(spare_reg_weight_19_15), .partial_sum_in(spare_reg_psum_19_15), .reg_activation(spare_reg_activation_20_15), .reg_weight(spare_reg_weight_20_15), .reg_partial_sum(spare_reg_psum_20_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_16( .activation_in(spare_reg_activation_20_15), .weight_in(spare_reg_weight_19_16), .partial_sum_in(spare_reg_psum_19_16), .reg_activation(spare_reg_activation_20_16), .reg_weight(spare_reg_weight_20_16), .reg_partial_sum(spare_reg_psum_20_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_17( .activation_in(spare_reg_activation_20_16), .weight_in(spare_reg_weight_19_17), .partial_sum_in(spare_reg_psum_19_17), .reg_activation(spare_reg_activation_20_17), .reg_weight(spare_reg_weight_20_17), .reg_partial_sum(spare_reg_psum_20_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_18( .activation_in(spare_reg_activation_20_17), .weight_in(spare_reg_weight_19_18), .partial_sum_in(spare_reg_psum_19_18), .reg_activation(spare_reg_activation_20_18), .reg_weight(spare_reg_weight_20_18), .reg_partial_sum(spare_reg_psum_20_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_19( .activation_in(spare_reg_activation_20_18), .weight_in(spare_reg_weight_19_19), .partial_sum_in(spare_reg_psum_19_19), .reg_activation(spare_reg_activation_20_19), .reg_weight(spare_reg_weight_20_19), .reg_partial_sum(spare_reg_psum_20_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_20( .activation_in(spare_reg_activation_20_19), .weight_in(spare_reg_weight_19_20), .partial_sum_in(spare_reg_psum_19_20), .reg_activation(spare_reg_activation_20_20), .reg_weight(spare_reg_weight_20_20), .reg_partial_sum(spare_reg_psum_20_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_21( .activation_in(spare_reg_activation_20_20), .weight_in(spare_reg_weight_19_21), .partial_sum_in(spare_reg_psum_19_21), .reg_activation(spare_reg_activation_20_21), .reg_weight(spare_reg_weight_20_21), .reg_partial_sum(spare_reg_psum_20_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_22( .activation_in(spare_reg_activation_20_21), .weight_in(spare_reg_weight_19_22), .partial_sum_in(spare_reg_psum_19_22), .reg_activation(spare_reg_activation_20_22), .reg_weight(spare_reg_weight_20_22), .reg_partial_sum(spare_reg_psum_20_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_23( .activation_in(spare_reg_activation_20_22), .weight_in(spare_reg_weight_19_23), .partial_sum_in(spare_reg_psum_19_23), .reg_activation(spare_reg_activation_20_23), .reg_weight(spare_reg_weight_20_23), .reg_partial_sum(spare_reg_psum_20_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_24( .activation_in(spare_reg_activation_20_23), .weight_in(spare_reg_weight_19_24), .partial_sum_in(spare_reg_psum_19_24), .reg_activation(spare_reg_activation_20_24), .reg_weight(spare_reg_weight_20_24), .reg_partial_sum(spare_reg_psum_20_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_25( .activation_in(spare_reg_activation_20_24), .weight_in(spare_reg_weight_19_25), .partial_sum_in(spare_reg_psum_19_25), .reg_activation(spare_reg_activation_20_25), .reg_weight(spare_reg_weight_20_25), .reg_partial_sum(spare_reg_psum_20_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_26( .activation_in(spare_reg_activation_20_25), .weight_in(spare_reg_weight_19_26), .partial_sum_in(spare_reg_psum_19_26), .reg_activation(spare_reg_activation_20_26), .reg_weight(spare_reg_weight_20_26), .reg_partial_sum(spare_reg_psum_20_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_27( .activation_in(spare_reg_activation_20_26), .weight_in(spare_reg_weight_19_27), .partial_sum_in(spare_reg_psum_19_27), .reg_activation(spare_reg_activation_20_27), .reg_weight(spare_reg_weight_20_27), .reg_partial_sum(spare_reg_psum_20_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_28( .activation_in(spare_reg_activation_20_27), .weight_in(spare_reg_weight_19_28), .partial_sum_in(spare_reg_psum_19_28), .reg_activation(spare_reg_activation_20_28), .reg_weight(spare_reg_weight_20_28), .reg_partial_sum(spare_reg_psum_20_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_29( .activation_in(spare_reg_activation_20_28), .weight_in(spare_reg_weight_19_29), .partial_sum_in(spare_reg_psum_19_29), .reg_activation(spare_reg_activation_20_29), .reg_weight(spare_reg_weight_20_29), .reg_partial_sum(spare_reg_psum_20_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_30( .activation_in(spare_reg_activation_20_29), .weight_in(spare_reg_weight_19_30), .partial_sum_in(spare_reg_psum_19_30), .reg_activation(spare_reg_activation_20_30), .reg_weight(spare_reg_weight_20_30), .reg_partial_sum(spare_reg_psum_20_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X20_31( .activation_in(spare_reg_activation_20_30), .weight_in(spare_reg_weight_19_31), .partial_sum_in(spare_reg_psum_19_31), .reg_weight(spare_reg_weight_20_31), .reg_partial_sum(spare_reg_psum_20_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_0( .activation_in(in_activation_21), .weight_in(spare_reg_weight_20_0), .partial_sum_in(spare_reg_psum_20_0), .reg_activation(spare_reg_activation_21_0), .reg_weight(spare_reg_weight_21_0), .reg_partial_sum(spare_reg_psum_21_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_1( .activation_in(spare_reg_activation_21_0), .weight_in(spare_reg_weight_20_1), .partial_sum_in(spare_reg_psum_20_1), .reg_activation(spare_reg_activation_21_1), .reg_weight(spare_reg_weight_21_1), .reg_partial_sum(spare_reg_psum_21_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_2( .activation_in(spare_reg_activation_21_1), .weight_in(spare_reg_weight_20_2), .partial_sum_in(spare_reg_psum_20_2), .reg_activation(spare_reg_activation_21_2), .reg_weight(spare_reg_weight_21_2), .reg_partial_sum(spare_reg_psum_21_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_3( .activation_in(spare_reg_activation_21_2), .weight_in(spare_reg_weight_20_3), .partial_sum_in(spare_reg_psum_20_3), .reg_activation(spare_reg_activation_21_3), .reg_weight(spare_reg_weight_21_3), .reg_partial_sum(spare_reg_psum_21_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_4( .activation_in(spare_reg_activation_21_3), .weight_in(spare_reg_weight_20_4), .partial_sum_in(spare_reg_psum_20_4), .reg_activation(spare_reg_activation_21_4), .reg_weight(spare_reg_weight_21_4), .reg_partial_sum(spare_reg_psum_21_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_5( .activation_in(spare_reg_activation_21_4), .weight_in(spare_reg_weight_20_5), .partial_sum_in(spare_reg_psum_20_5), .reg_activation(spare_reg_activation_21_5), .reg_weight(spare_reg_weight_21_5), .reg_partial_sum(spare_reg_psum_21_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_6( .activation_in(spare_reg_activation_21_5), .weight_in(spare_reg_weight_20_6), .partial_sum_in(spare_reg_psum_20_6), .reg_activation(spare_reg_activation_21_6), .reg_weight(spare_reg_weight_21_6), .reg_partial_sum(spare_reg_psum_21_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_7( .activation_in(spare_reg_activation_21_6), .weight_in(spare_reg_weight_20_7), .partial_sum_in(spare_reg_psum_20_7), .reg_activation(spare_reg_activation_21_7), .reg_weight(spare_reg_weight_21_7), .reg_partial_sum(spare_reg_psum_21_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_8( .activation_in(spare_reg_activation_21_7), .weight_in(spare_reg_weight_20_8), .partial_sum_in(spare_reg_psum_20_8), .reg_activation(spare_reg_activation_21_8), .reg_weight(spare_reg_weight_21_8), .reg_partial_sum(spare_reg_psum_21_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_9( .activation_in(spare_reg_activation_21_8), .weight_in(spare_reg_weight_20_9), .partial_sum_in(spare_reg_psum_20_9), .reg_activation(spare_reg_activation_21_9), .reg_weight(spare_reg_weight_21_9), .reg_partial_sum(spare_reg_psum_21_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_10( .activation_in(spare_reg_activation_21_9), .weight_in(spare_reg_weight_20_10), .partial_sum_in(spare_reg_psum_20_10), .reg_activation(spare_reg_activation_21_10), .reg_weight(spare_reg_weight_21_10), .reg_partial_sum(spare_reg_psum_21_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_11( .activation_in(spare_reg_activation_21_10), .weight_in(spare_reg_weight_20_11), .partial_sum_in(spare_reg_psum_20_11), .reg_activation(spare_reg_activation_21_11), .reg_weight(spare_reg_weight_21_11), .reg_partial_sum(spare_reg_psum_21_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_12( .activation_in(spare_reg_activation_21_11), .weight_in(spare_reg_weight_20_12), .partial_sum_in(spare_reg_psum_20_12), .reg_activation(spare_reg_activation_21_12), .reg_weight(spare_reg_weight_21_12), .reg_partial_sum(spare_reg_psum_21_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_13( .activation_in(spare_reg_activation_21_12), .weight_in(spare_reg_weight_20_13), .partial_sum_in(spare_reg_psum_20_13), .reg_activation(spare_reg_activation_21_13), .reg_weight(spare_reg_weight_21_13), .reg_partial_sum(spare_reg_psum_21_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_14( .activation_in(spare_reg_activation_21_13), .weight_in(spare_reg_weight_20_14), .partial_sum_in(spare_reg_psum_20_14), .reg_activation(spare_reg_activation_21_14), .reg_weight(spare_reg_weight_21_14), .reg_partial_sum(spare_reg_psum_21_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_15( .activation_in(spare_reg_activation_21_14), .weight_in(spare_reg_weight_20_15), .partial_sum_in(spare_reg_psum_20_15), .reg_activation(spare_reg_activation_21_15), .reg_weight(spare_reg_weight_21_15), .reg_partial_sum(spare_reg_psum_21_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_16( .activation_in(spare_reg_activation_21_15), .weight_in(spare_reg_weight_20_16), .partial_sum_in(spare_reg_psum_20_16), .reg_activation(spare_reg_activation_21_16), .reg_weight(spare_reg_weight_21_16), .reg_partial_sum(spare_reg_psum_21_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_17( .activation_in(spare_reg_activation_21_16), .weight_in(spare_reg_weight_20_17), .partial_sum_in(spare_reg_psum_20_17), .reg_activation(spare_reg_activation_21_17), .reg_weight(spare_reg_weight_21_17), .reg_partial_sum(spare_reg_psum_21_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_18( .activation_in(spare_reg_activation_21_17), .weight_in(spare_reg_weight_20_18), .partial_sum_in(spare_reg_psum_20_18), .reg_activation(spare_reg_activation_21_18), .reg_weight(spare_reg_weight_21_18), .reg_partial_sum(spare_reg_psum_21_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_19( .activation_in(spare_reg_activation_21_18), .weight_in(spare_reg_weight_20_19), .partial_sum_in(spare_reg_psum_20_19), .reg_activation(spare_reg_activation_21_19), .reg_weight(spare_reg_weight_21_19), .reg_partial_sum(spare_reg_psum_21_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_20( .activation_in(spare_reg_activation_21_19), .weight_in(spare_reg_weight_20_20), .partial_sum_in(spare_reg_psum_20_20), .reg_activation(spare_reg_activation_21_20), .reg_weight(spare_reg_weight_21_20), .reg_partial_sum(spare_reg_psum_21_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_21( .activation_in(spare_reg_activation_21_20), .weight_in(spare_reg_weight_20_21), .partial_sum_in(spare_reg_psum_20_21), .reg_activation(spare_reg_activation_21_21), .reg_weight(spare_reg_weight_21_21), .reg_partial_sum(spare_reg_psum_21_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_22( .activation_in(spare_reg_activation_21_21), .weight_in(spare_reg_weight_20_22), .partial_sum_in(spare_reg_psum_20_22), .reg_activation(spare_reg_activation_21_22), .reg_weight(spare_reg_weight_21_22), .reg_partial_sum(spare_reg_psum_21_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_23( .activation_in(spare_reg_activation_21_22), .weight_in(spare_reg_weight_20_23), .partial_sum_in(spare_reg_psum_20_23), .reg_activation(spare_reg_activation_21_23), .reg_weight(spare_reg_weight_21_23), .reg_partial_sum(spare_reg_psum_21_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_24( .activation_in(spare_reg_activation_21_23), .weight_in(spare_reg_weight_20_24), .partial_sum_in(spare_reg_psum_20_24), .reg_activation(spare_reg_activation_21_24), .reg_weight(spare_reg_weight_21_24), .reg_partial_sum(spare_reg_psum_21_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_25( .activation_in(spare_reg_activation_21_24), .weight_in(spare_reg_weight_20_25), .partial_sum_in(spare_reg_psum_20_25), .reg_activation(spare_reg_activation_21_25), .reg_weight(spare_reg_weight_21_25), .reg_partial_sum(spare_reg_psum_21_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_26( .activation_in(spare_reg_activation_21_25), .weight_in(spare_reg_weight_20_26), .partial_sum_in(spare_reg_psum_20_26), .reg_activation(spare_reg_activation_21_26), .reg_weight(spare_reg_weight_21_26), .reg_partial_sum(spare_reg_psum_21_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_27( .activation_in(spare_reg_activation_21_26), .weight_in(spare_reg_weight_20_27), .partial_sum_in(spare_reg_psum_20_27), .reg_activation(spare_reg_activation_21_27), .reg_weight(spare_reg_weight_21_27), .reg_partial_sum(spare_reg_psum_21_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_28( .activation_in(spare_reg_activation_21_27), .weight_in(spare_reg_weight_20_28), .partial_sum_in(spare_reg_psum_20_28), .reg_activation(spare_reg_activation_21_28), .reg_weight(spare_reg_weight_21_28), .reg_partial_sum(spare_reg_psum_21_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_29( .activation_in(spare_reg_activation_21_28), .weight_in(spare_reg_weight_20_29), .partial_sum_in(spare_reg_psum_20_29), .reg_activation(spare_reg_activation_21_29), .reg_weight(spare_reg_weight_21_29), .reg_partial_sum(spare_reg_psum_21_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_30( .activation_in(spare_reg_activation_21_29), .weight_in(spare_reg_weight_20_30), .partial_sum_in(spare_reg_psum_20_30), .reg_activation(spare_reg_activation_21_30), .reg_weight(spare_reg_weight_21_30), .reg_partial_sum(spare_reg_psum_21_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X21_31( .activation_in(spare_reg_activation_21_30), .weight_in(spare_reg_weight_20_31), .partial_sum_in(spare_reg_psum_20_31), .reg_weight(spare_reg_weight_21_31), .reg_partial_sum(spare_reg_psum_21_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_0( .activation_in(in_activation_22), .weight_in(spare_reg_weight_21_0), .partial_sum_in(spare_reg_psum_21_0), .reg_activation(spare_reg_activation_22_0), .reg_weight(spare_reg_weight_22_0), .reg_partial_sum(spare_reg_psum_22_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_1( .activation_in(spare_reg_activation_22_0), .weight_in(spare_reg_weight_21_1), .partial_sum_in(spare_reg_psum_21_1), .reg_activation(spare_reg_activation_22_1), .reg_weight(spare_reg_weight_22_1), .reg_partial_sum(spare_reg_psum_22_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_2( .activation_in(spare_reg_activation_22_1), .weight_in(spare_reg_weight_21_2), .partial_sum_in(spare_reg_psum_21_2), .reg_activation(spare_reg_activation_22_2), .reg_weight(spare_reg_weight_22_2), .reg_partial_sum(spare_reg_psum_22_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_3( .activation_in(spare_reg_activation_22_2), .weight_in(spare_reg_weight_21_3), .partial_sum_in(spare_reg_psum_21_3), .reg_activation(spare_reg_activation_22_3), .reg_weight(spare_reg_weight_22_3), .reg_partial_sum(spare_reg_psum_22_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_4( .activation_in(spare_reg_activation_22_3), .weight_in(spare_reg_weight_21_4), .partial_sum_in(spare_reg_psum_21_4), .reg_activation(spare_reg_activation_22_4), .reg_weight(spare_reg_weight_22_4), .reg_partial_sum(spare_reg_psum_22_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_5( .activation_in(spare_reg_activation_22_4), .weight_in(spare_reg_weight_21_5), .partial_sum_in(spare_reg_psum_21_5), .reg_activation(spare_reg_activation_22_5), .reg_weight(spare_reg_weight_22_5), .reg_partial_sum(spare_reg_psum_22_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_6( .activation_in(spare_reg_activation_22_5), .weight_in(spare_reg_weight_21_6), .partial_sum_in(spare_reg_psum_21_6), .reg_activation(spare_reg_activation_22_6), .reg_weight(spare_reg_weight_22_6), .reg_partial_sum(spare_reg_psum_22_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_7( .activation_in(spare_reg_activation_22_6), .weight_in(spare_reg_weight_21_7), .partial_sum_in(spare_reg_psum_21_7), .reg_activation(spare_reg_activation_22_7), .reg_weight(spare_reg_weight_22_7), .reg_partial_sum(spare_reg_psum_22_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_8( .activation_in(spare_reg_activation_22_7), .weight_in(spare_reg_weight_21_8), .partial_sum_in(spare_reg_psum_21_8), .reg_activation(spare_reg_activation_22_8), .reg_weight(spare_reg_weight_22_8), .reg_partial_sum(spare_reg_psum_22_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_9( .activation_in(spare_reg_activation_22_8), .weight_in(spare_reg_weight_21_9), .partial_sum_in(spare_reg_psum_21_9), .reg_activation(spare_reg_activation_22_9), .reg_weight(spare_reg_weight_22_9), .reg_partial_sum(spare_reg_psum_22_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_10( .activation_in(spare_reg_activation_22_9), .weight_in(spare_reg_weight_21_10), .partial_sum_in(spare_reg_psum_21_10), .reg_activation(spare_reg_activation_22_10), .reg_weight(spare_reg_weight_22_10), .reg_partial_sum(spare_reg_psum_22_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_11( .activation_in(spare_reg_activation_22_10), .weight_in(spare_reg_weight_21_11), .partial_sum_in(spare_reg_psum_21_11), .reg_activation(spare_reg_activation_22_11), .reg_weight(spare_reg_weight_22_11), .reg_partial_sum(spare_reg_psum_22_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_12( .activation_in(spare_reg_activation_22_11), .weight_in(spare_reg_weight_21_12), .partial_sum_in(spare_reg_psum_21_12), .reg_activation(spare_reg_activation_22_12), .reg_weight(spare_reg_weight_22_12), .reg_partial_sum(spare_reg_psum_22_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_13( .activation_in(spare_reg_activation_22_12), .weight_in(spare_reg_weight_21_13), .partial_sum_in(spare_reg_psum_21_13), .reg_activation(spare_reg_activation_22_13), .reg_weight(spare_reg_weight_22_13), .reg_partial_sum(spare_reg_psum_22_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_14( .activation_in(spare_reg_activation_22_13), .weight_in(spare_reg_weight_21_14), .partial_sum_in(spare_reg_psum_21_14), .reg_activation(spare_reg_activation_22_14), .reg_weight(spare_reg_weight_22_14), .reg_partial_sum(spare_reg_psum_22_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_15( .activation_in(spare_reg_activation_22_14), .weight_in(spare_reg_weight_21_15), .partial_sum_in(spare_reg_psum_21_15), .reg_activation(spare_reg_activation_22_15), .reg_weight(spare_reg_weight_22_15), .reg_partial_sum(spare_reg_psum_22_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_16( .activation_in(spare_reg_activation_22_15), .weight_in(spare_reg_weight_21_16), .partial_sum_in(spare_reg_psum_21_16), .reg_activation(spare_reg_activation_22_16), .reg_weight(spare_reg_weight_22_16), .reg_partial_sum(spare_reg_psum_22_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_17( .activation_in(spare_reg_activation_22_16), .weight_in(spare_reg_weight_21_17), .partial_sum_in(spare_reg_psum_21_17), .reg_activation(spare_reg_activation_22_17), .reg_weight(spare_reg_weight_22_17), .reg_partial_sum(spare_reg_psum_22_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_18( .activation_in(spare_reg_activation_22_17), .weight_in(spare_reg_weight_21_18), .partial_sum_in(spare_reg_psum_21_18), .reg_activation(spare_reg_activation_22_18), .reg_weight(spare_reg_weight_22_18), .reg_partial_sum(spare_reg_psum_22_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_19( .activation_in(spare_reg_activation_22_18), .weight_in(spare_reg_weight_21_19), .partial_sum_in(spare_reg_psum_21_19), .reg_activation(spare_reg_activation_22_19), .reg_weight(spare_reg_weight_22_19), .reg_partial_sum(spare_reg_psum_22_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_20( .activation_in(spare_reg_activation_22_19), .weight_in(spare_reg_weight_21_20), .partial_sum_in(spare_reg_psum_21_20), .reg_activation(spare_reg_activation_22_20), .reg_weight(spare_reg_weight_22_20), .reg_partial_sum(spare_reg_psum_22_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_21( .activation_in(spare_reg_activation_22_20), .weight_in(spare_reg_weight_21_21), .partial_sum_in(spare_reg_psum_21_21), .reg_activation(spare_reg_activation_22_21), .reg_weight(spare_reg_weight_22_21), .reg_partial_sum(spare_reg_psum_22_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_22( .activation_in(spare_reg_activation_22_21), .weight_in(spare_reg_weight_21_22), .partial_sum_in(spare_reg_psum_21_22), .reg_activation(spare_reg_activation_22_22), .reg_weight(spare_reg_weight_22_22), .reg_partial_sum(spare_reg_psum_22_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_23( .activation_in(spare_reg_activation_22_22), .weight_in(spare_reg_weight_21_23), .partial_sum_in(spare_reg_psum_21_23), .reg_activation(spare_reg_activation_22_23), .reg_weight(spare_reg_weight_22_23), .reg_partial_sum(spare_reg_psum_22_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_24( .activation_in(spare_reg_activation_22_23), .weight_in(spare_reg_weight_21_24), .partial_sum_in(spare_reg_psum_21_24), .reg_activation(spare_reg_activation_22_24), .reg_weight(spare_reg_weight_22_24), .reg_partial_sum(spare_reg_psum_22_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_25( .activation_in(spare_reg_activation_22_24), .weight_in(spare_reg_weight_21_25), .partial_sum_in(spare_reg_psum_21_25), .reg_activation(spare_reg_activation_22_25), .reg_weight(spare_reg_weight_22_25), .reg_partial_sum(spare_reg_psum_22_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_26( .activation_in(spare_reg_activation_22_25), .weight_in(spare_reg_weight_21_26), .partial_sum_in(spare_reg_psum_21_26), .reg_activation(spare_reg_activation_22_26), .reg_weight(spare_reg_weight_22_26), .reg_partial_sum(spare_reg_psum_22_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_27( .activation_in(spare_reg_activation_22_26), .weight_in(spare_reg_weight_21_27), .partial_sum_in(spare_reg_psum_21_27), .reg_activation(spare_reg_activation_22_27), .reg_weight(spare_reg_weight_22_27), .reg_partial_sum(spare_reg_psum_22_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_28( .activation_in(spare_reg_activation_22_27), .weight_in(spare_reg_weight_21_28), .partial_sum_in(spare_reg_psum_21_28), .reg_activation(spare_reg_activation_22_28), .reg_weight(spare_reg_weight_22_28), .reg_partial_sum(spare_reg_psum_22_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_29( .activation_in(spare_reg_activation_22_28), .weight_in(spare_reg_weight_21_29), .partial_sum_in(spare_reg_psum_21_29), .reg_activation(spare_reg_activation_22_29), .reg_weight(spare_reg_weight_22_29), .reg_partial_sum(spare_reg_psum_22_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_30( .activation_in(spare_reg_activation_22_29), .weight_in(spare_reg_weight_21_30), .partial_sum_in(spare_reg_psum_21_30), .reg_activation(spare_reg_activation_22_30), .reg_weight(spare_reg_weight_22_30), .reg_partial_sum(spare_reg_psum_22_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X22_31( .activation_in(spare_reg_activation_22_30), .weight_in(spare_reg_weight_21_31), .partial_sum_in(spare_reg_psum_21_31), .reg_weight(spare_reg_weight_22_31), .reg_partial_sum(spare_reg_psum_22_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_0( .activation_in(in_activation_23), .weight_in(spare_reg_weight_22_0), .partial_sum_in(spare_reg_psum_22_0), .reg_activation(spare_reg_activation_23_0), .reg_weight(spare_reg_weight_23_0), .reg_partial_sum(spare_reg_psum_23_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_1( .activation_in(spare_reg_activation_23_0), .weight_in(spare_reg_weight_22_1), .partial_sum_in(spare_reg_psum_22_1), .reg_activation(spare_reg_activation_23_1), .reg_weight(spare_reg_weight_23_1), .reg_partial_sum(spare_reg_psum_23_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_2( .activation_in(spare_reg_activation_23_1), .weight_in(spare_reg_weight_22_2), .partial_sum_in(spare_reg_psum_22_2), .reg_activation(spare_reg_activation_23_2), .reg_weight(spare_reg_weight_23_2), .reg_partial_sum(spare_reg_psum_23_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_3( .activation_in(spare_reg_activation_23_2), .weight_in(spare_reg_weight_22_3), .partial_sum_in(spare_reg_psum_22_3), .reg_activation(spare_reg_activation_23_3), .reg_weight(spare_reg_weight_23_3), .reg_partial_sum(spare_reg_psum_23_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_4( .activation_in(spare_reg_activation_23_3), .weight_in(spare_reg_weight_22_4), .partial_sum_in(spare_reg_psum_22_4), .reg_activation(spare_reg_activation_23_4), .reg_weight(spare_reg_weight_23_4), .reg_partial_sum(spare_reg_psum_23_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_5( .activation_in(spare_reg_activation_23_4), .weight_in(spare_reg_weight_22_5), .partial_sum_in(spare_reg_psum_22_5), .reg_activation(spare_reg_activation_23_5), .reg_weight(spare_reg_weight_23_5), .reg_partial_sum(spare_reg_psum_23_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_6( .activation_in(spare_reg_activation_23_5), .weight_in(spare_reg_weight_22_6), .partial_sum_in(spare_reg_psum_22_6), .reg_activation(spare_reg_activation_23_6), .reg_weight(spare_reg_weight_23_6), .reg_partial_sum(spare_reg_psum_23_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_7( .activation_in(spare_reg_activation_23_6), .weight_in(spare_reg_weight_22_7), .partial_sum_in(spare_reg_psum_22_7), .reg_activation(spare_reg_activation_23_7), .reg_weight(spare_reg_weight_23_7), .reg_partial_sum(spare_reg_psum_23_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_8( .activation_in(spare_reg_activation_23_7), .weight_in(spare_reg_weight_22_8), .partial_sum_in(spare_reg_psum_22_8), .reg_activation(spare_reg_activation_23_8), .reg_weight(spare_reg_weight_23_8), .reg_partial_sum(spare_reg_psum_23_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_9( .activation_in(spare_reg_activation_23_8), .weight_in(spare_reg_weight_22_9), .partial_sum_in(spare_reg_psum_22_9), .reg_activation(spare_reg_activation_23_9), .reg_weight(spare_reg_weight_23_9), .reg_partial_sum(spare_reg_psum_23_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_10( .activation_in(spare_reg_activation_23_9), .weight_in(spare_reg_weight_22_10), .partial_sum_in(spare_reg_psum_22_10), .reg_activation(spare_reg_activation_23_10), .reg_weight(spare_reg_weight_23_10), .reg_partial_sum(spare_reg_psum_23_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_11( .activation_in(spare_reg_activation_23_10), .weight_in(spare_reg_weight_22_11), .partial_sum_in(spare_reg_psum_22_11), .reg_activation(spare_reg_activation_23_11), .reg_weight(spare_reg_weight_23_11), .reg_partial_sum(spare_reg_psum_23_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_12( .activation_in(spare_reg_activation_23_11), .weight_in(spare_reg_weight_22_12), .partial_sum_in(spare_reg_psum_22_12), .reg_activation(spare_reg_activation_23_12), .reg_weight(spare_reg_weight_23_12), .reg_partial_sum(spare_reg_psum_23_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_13( .activation_in(spare_reg_activation_23_12), .weight_in(spare_reg_weight_22_13), .partial_sum_in(spare_reg_psum_22_13), .reg_activation(spare_reg_activation_23_13), .reg_weight(spare_reg_weight_23_13), .reg_partial_sum(spare_reg_psum_23_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_14( .activation_in(spare_reg_activation_23_13), .weight_in(spare_reg_weight_22_14), .partial_sum_in(spare_reg_psum_22_14), .reg_activation(spare_reg_activation_23_14), .reg_weight(spare_reg_weight_23_14), .reg_partial_sum(spare_reg_psum_23_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_15( .activation_in(spare_reg_activation_23_14), .weight_in(spare_reg_weight_22_15), .partial_sum_in(spare_reg_psum_22_15), .reg_activation(spare_reg_activation_23_15), .reg_weight(spare_reg_weight_23_15), .reg_partial_sum(spare_reg_psum_23_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_16( .activation_in(spare_reg_activation_23_15), .weight_in(spare_reg_weight_22_16), .partial_sum_in(spare_reg_psum_22_16), .reg_activation(spare_reg_activation_23_16), .reg_weight(spare_reg_weight_23_16), .reg_partial_sum(spare_reg_psum_23_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_17( .activation_in(spare_reg_activation_23_16), .weight_in(spare_reg_weight_22_17), .partial_sum_in(spare_reg_psum_22_17), .reg_activation(spare_reg_activation_23_17), .reg_weight(spare_reg_weight_23_17), .reg_partial_sum(spare_reg_psum_23_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_18( .activation_in(spare_reg_activation_23_17), .weight_in(spare_reg_weight_22_18), .partial_sum_in(spare_reg_psum_22_18), .reg_activation(spare_reg_activation_23_18), .reg_weight(spare_reg_weight_23_18), .reg_partial_sum(spare_reg_psum_23_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_19( .activation_in(spare_reg_activation_23_18), .weight_in(spare_reg_weight_22_19), .partial_sum_in(spare_reg_psum_22_19), .reg_activation(spare_reg_activation_23_19), .reg_weight(spare_reg_weight_23_19), .reg_partial_sum(spare_reg_psum_23_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_20( .activation_in(spare_reg_activation_23_19), .weight_in(spare_reg_weight_22_20), .partial_sum_in(spare_reg_psum_22_20), .reg_activation(spare_reg_activation_23_20), .reg_weight(spare_reg_weight_23_20), .reg_partial_sum(spare_reg_psum_23_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_21( .activation_in(spare_reg_activation_23_20), .weight_in(spare_reg_weight_22_21), .partial_sum_in(spare_reg_psum_22_21), .reg_activation(spare_reg_activation_23_21), .reg_weight(spare_reg_weight_23_21), .reg_partial_sum(spare_reg_psum_23_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_22( .activation_in(spare_reg_activation_23_21), .weight_in(spare_reg_weight_22_22), .partial_sum_in(spare_reg_psum_22_22), .reg_activation(spare_reg_activation_23_22), .reg_weight(spare_reg_weight_23_22), .reg_partial_sum(spare_reg_psum_23_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_23( .activation_in(spare_reg_activation_23_22), .weight_in(spare_reg_weight_22_23), .partial_sum_in(spare_reg_psum_22_23), .reg_activation(spare_reg_activation_23_23), .reg_weight(spare_reg_weight_23_23), .reg_partial_sum(spare_reg_psum_23_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_24( .activation_in(spare_reg_activation_23_23), .weight_in(spare_reg_weight_22_24), .partial_sum_in(spare_reg_psum_22_24), .reg_activation(spare_reg_activation_23_24), .reg_weight(spare_reg_weight_23_24), .reg_partial_sum(spare_reg_psum_23_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_25( .activation_in(spare_reg_activation_23_24), .weight_in(spare_reg_weight_22_25), .partial_sum_in(spare_reg_psum_22_25), .reg_activation(spare_reg_activation_23_25), .reg_weight(spare_reg_weight_23_25), .reg_partial_sum(spare_reg_psum_23_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_26( .activation_in(spare_reg_activation_23_25), .weight_in(spare_reg_weight_22_26), .partial_sum_in(spare_reg_psum_22_26), .reg_activation(spare_reg_activation_23_26), .reg_weight(spare_reg_weight_23_26), .reg_partial_sum(spare_reg_psum_23_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_27( .activation_in(spare_reg_activation_23_26), .weight_in(spare_reg_weight_22_27), .partial_sum_in(spare_reg_psum_22_27), .reg_activation(spare_reg_activation_23_27), .reg_weight(spare_reg_weight_23_27), .reg_partial_sum(spare_reg_psum_23_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_28( .activation_in(spare_reg_activation_23_27), .weight_in(spare_reg_weight_22_28), .partial_sum_in(spare_reg_psum_22_28), .reg_activation(spare_reg_activation_23_28), .reg_weight(spare_reg_weight_23_28), .reg_partial_sum(spare_reg_psum_23_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_29( .activation_in(spare_reg_activation_23_28), .weight_in(spare_reg_weight_22_29), .partial_sum_in(spare_reg_psum_22_29), .reg_activation(spare_reg_activation_23_29), .reg_weight(spare_reg_weight_23_29), .reg_partial_sum(spare_reg_psum_23_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_30( .activation_in(spare_reg_activation_23_29), .weight_in(spare_reg_weight_22_30), .partial_sum_in(spare_reg_psum_22_30), .reg_activation(spare_reg_activation_23_30), .reg_weight(spare_reg_weight_23_30), .reg_partial_sum(spare_reg_psum_23_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X23_31( .activation_in(spare_reg_activation_23_30), .weight_in(spare_reg_weight_22_31), .partial_sum_in(spare_reg_psum_22_31), .reg_weight(spare_reg_weight_23_31), .reg_partial_sum(spare_reg_psum_23_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_0( .activation_in(in_activation_24), .weight_in(spare_reg_weight_23_0), .partial_sum_in(spare_reg_psum_23_0), .reg_activation(spare_reg_activation_24_0), .reg_weight(spare_reg_weight_24_0), .reg_partial_sum(spare_reg_psum_24_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_1( .activation_in(spare_reg_activation_24_0), .weight_in(spare_reg_weight_23_1), .partial_sum_in(spare_reg_psum_23_1), .reg_activation(spare_reg_activation_24_1), .reg_weight(spare_reg_weight_24_1), .reg_partial_sum(spare_reg_psum_24_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_2( .activation_in(spare_reg_activation_24_1), .weight_in(spare_reg_weight_23_2), .partial_sum_in(spare_reg_psum_23_2), .reg_activation(spare_reg_activation_24_2), .reg_weight(spare_reg_weight_24_2), .reg_partial_sum(spare_reg_psum_24_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_3( .activation_in(spare_reg_activation_24_2), .weight_in(spare_reg_weight_23_3), .partial_sum_in(spare_reg_psum_23_3), .reg_activation(spare_reg_activation_24_3), .reg_weight(spare_reg_weight_24_3), .reg_partial_sum(spare_reg_psum_24_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_4( .activation_in(spare_reg_activation_24_3), .weight_in(spare_reg_weight_23_4), .partial_sum_in(spare_reg_psum_23_4), .reg_activation(spare_reg_activation_24_4), .reg_weight(spare_reg_weight_24_4), .reg_partial_sum(spare_reg_psum_24_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_5( .activation_in(spare_reg_activation_24_4), .weight_in(spare_reg_weight_23_5), .partial_sum_in(spare_reg_psum_23_5), .reg_activation(spare_reg_activation_24_5), .reg_weight(spare_reg_weight_24_5), .reg_partial_sum(spare_reg_psum_24_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_6( .activation_in(spare_reg_activation_24_5), .weight_in(spare_reg_weight_23_6), .partial_sum_in(spare_reg_psum_23_6), .reg_activation(spare_reg_activation_24_6), .reg_weight(spare_reg_weight_24_6), .reg_partial_sum(spare_reg_psum_24_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_7( .activation_in(spare_reg_activation_24_6), .weight_in(spare_reg_weight_23_7), .partial_sum_in(spare_reg_psum_23_7), .reg_activation(spare_reg_activation_24_7), .reg_weight(spare_reg_weight_24_7), .reg_partial_sum(spare_reg_psum_24_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_8( .activation_in(spare_reg_activation_24_7), .weight_in(spare_reg_weight_23_8), .partial_sum_in(spare_reg_psum_23_8), .reg_activation(spare_reg_activation_24_8), .reg_weight(spare_reg_weight_24_8), .reg_partial_sum(spare_reg_psum_24_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_9( .activation_in(spare_reg_activation_24_8), .weight_in(spare_reg_weight_23_9), .partial_sum_in(spare_reg_psum_23_9), .reg_activation(spare_reg_activation_24_9), .reg_weight(spare_reg_weight_24_9), .reg_partial_sum(spare_reg_psum_24_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_10( .activation_in(spare_reg_activation_24_9), .weight_in(spare_reg_weight_23_10), .partial_sum_in(spare_reg_psum_23_10), .reg_activation(spare_reg_activation_24_10), .reg_weight(spare_reg_weight_24_10), .reg_partial_sum(spare_reg_psum_24_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_11( .activation_in(spare_reg_activation_24_10), .weight_in(spare_reg_weight_23_11), .partial_sum_in(spare_reg_psum_23_11), .reg_activation(spare_reg_activation_24_11), .reg_weight(spare_reg_weight_24_11), .reg_partial_sum(spare_reg_psum_24_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_12( .activation_in(spare_reg_activation_24_11), .weight_in(spare_reg_weight_23_12), .partial_sum_in(spare_reg_psum_23_12), .reg_activation(spare_reg_activation_24_12), .reg_weight(spare_reg_weight_24_12), .reg_partial_sum(spare_reg_psum_24_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_13( .activation_in(spare_reg_activation_24_12), .weight_in(spare_reg_weight_23_13), .partial_sum_in(spare_reg_psum_23_13), .reg_activation(spare_reg_activation_24_13), .reg_weight(spare_reg_weight_24_13), .reg_partial_sum(spare_reg_psum_24_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_14( .activation_in(spare_reg_activation_24_13), .weight_in(spare_reg_weight_23_14), .partial_sum_in(spare_reg_psum_23_14), .reg_activation(spare_reg_activation_24_14), .reg_weight(spare_reg_weight_24_14), .reg_partial_sum(spare_reg_psum_24_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_15( .activation_in(spare_reg_activation_24_14), .weight_in(spare_reg_weight_23_15), .partial_sum_in(spare_reg_psum_23_15), .reg_activation(spare_reg_activation_24_15), .reg_weight(spare_reg_weight_24_15), .reg_partial_sum(spare_reg_psum_24_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_16( .activation_in(spare_reg_activation_24_15), .weight_in(spare_reg_weight_23_16), .partial_sum_in(spare_reg_psum_23_16), .reg_activation(spare_reg_activation_24_16), .reg_weight(spare_reg_weight_24_16), .reg_partial_sum(spare_reg_psum_24_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_17( .activation_in(spare_reg_activation_24_16), .weight_in(spare_reg_weight_23_17), .partial_sum_in(spare_reg_psum_23_17), .reg_activation(spare_reg_activation_24_17), .reg_weight(spare_reg_weight_24_17), .reg_partial_sum(spare_reg_psum_24_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_18( .activation_in(spare_reg_activation_24_17), .weight_in(spare_reg_weight_23_18), .partial_sum_in(spare_reg_psum_23_18), .reg_activation(spare_reg_activation_24_18), .reg_weight(spare_reg_weight_24_18), .reg_partial_sum(spare_reg_psum_24_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_19( .activation_in(spare_reg_activation_24_18), .weight_in(spare_reg_weight_23_19), .partial_sum_in(spare_reg_psum_23_19), .reg_activation(spare_reg_activation_24_19), .reg_weight(spare_reg_weight_24_19), .reg_partial_sum(spare_reg_psum_24_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_20( .activation_in(spare_reg_activation_24_19), .weight_in(spare_reg_weight_23_20), .partial_sum_in(spare_reg_psum_23_20), .reg_activation(spare_reg_activation_24_20), .reg_weight(spare_reg_weight_24_20), .reg_partial_sum(spare_reg_psum_24_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_21( .activation_in(spare_reg_activation_24_20), .weight_in(spare_reg_weight_23_21), .partial_sum_in(spare_reg_psum_23_21), .reg_activation(spare_reg_activation_24_21), .reg_weight(spare_reg_weight_24_21), .reg_partial_sum(spare_reg_psum_24_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_22( .activation_in(spare_reg_activation_24_21), .weight_in(spare_reg_weight_23_22), .partial_sum_in(spare_reg_psum_23_22), .reg_activation(spare_reg_activation_24_22), .reg_weight(spare_reg_weight_24_22), .reg_partial_sum(spare_reg_psum_24_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_23( .activation_in(spare_reg_activation_24_22), .weight_in(spare_reg_weight_23_23), .partial_sum_in(spare_reg_psum_23_23), .reg_activation(spare_reg_activation_24_23), .reg_weight(spare_reg_weight_24_23), .reg_partial_sum(spare_reg_psum_24_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_24( .activation_in(spare_reg_activation_24_23), .weight_in(spare_reg_weight_23_24), .partial_sum_in(spare_reg_psum_23_24), .reg_activation(spare_reg_activation_24_24), .reg_weight(spare_reg_weight_24_24), .reg_partial_sum(spare_reg_psum_24_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_25( .activation_in(spare_reg_activation_24_24), .weight_in(spare_reg_weight_23_25), .partial_sum_in(spare_reg_psum_23_25), .reg_activation(spare_reg_activation_24_25), .reg_weight(spare_reg_weight_24_25), .reg_partial_sum(spare_reg_psum_24_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_26( .activation_in(spare_reg_activation_24_25), .weight_in(spare_reg_weight_23_26), .partial_sum_in(spare_reg_psum_23_26), .reg_activation(spare_reg_activation_24_26), .reg_weight(spare_reg_weight_24_26), .reg_partial_sum(spare_reg_psum_24_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_27( .activation_in(spare_reg_activation_24_26), .weight_in(spare_reg_weight_23_27), .partial_sum_in(spare_reg_psum_23_27), .reg_activation(spare_reg_activation_24_27), .reg_weight(spare_reg_weight_24_27), .reg_partial_sum(spare_reg_psum_24_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_28( .activation_in(spare_reg_activation_24_27), .weight_in(spare_reg_weight_23_28), .partial_sum_in(spare_reg_psum_23_28), .reg_activation(spare_reg_activation_24_28), .reg_weight(spare_reg_weight_24_28), .reg_partial_sum(spare_reg_psum_24_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_29( .activation_in(spare_reg_activation_24_28), .weight_in(spare_reg_weight_23_29), .partial_sum_in(spare_reg_psum_23_29), .reg_activation(spare_reg_activation_24_29), .reg_weight(spare_reg_weight_24_29), .reg_partial_sum(spare_reg_psum_24_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_30( .activation_in(spare_reg_activation_24_29), .weight_in(spare_reg_weight_23_30), .partial_sum_in(spare_reg_psum_23_30), .reg_activation(spare_reg_activation_24_30), .reg_weight(spare_reg_weight_24_30), .reg_partial_sum(spare_reg_psum_24_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X24_31( .activation_in(spare_reg_activation_24_30), .weight_in(spare_reg_weight_23_31), .partial_sum_in(spare_reg_psum_23_31), .reg_weight(spare_reg_weight_24_31), .reg_partial_sum(spare_reg_psum_24_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_0( .activation_in(in_activation_25), .weight_in(spare_reg_weight_24_0), .partial_sum_in(spare_reg_psum_24_0), .reg_activation(spare_reg_activation_25_0), .reg_weight(spare_reg_weight_25_0), .reg_partial_sum(spare_reg_psum_25_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_1( .activation_in(spare_reg_activation_25_0), .weight_in(spare_reg_weight_24_1), .partial_sum_in(spare_reg_psum_24_1), .reg_activation(spare_reg_activation_25_1), .reg_weight(spare_reg_weight_25_1), .reg_partial_sum(spare_reg_psum_25_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_2( .activation_in(spare_reg_activation_25_1), .weight_in(spare_reg_weight_24_2), .partial_sum_in(spare_reg_psum_24_2), .reg_activation(spare_reg_activation_25_2), .reg_weight(spare_reg_weight_25_2), .reg_partial_sum(spare_reg_psum_25_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_3( .activation_in(spare_reg_activation_25_2), .weight_in(spare_reg_weight_24_3), .partial_sum_in(spare_reg_psum_24_3), .reg_activation(spare_reg_activation_25_3), .reg_weight(spare_reg_weight_25_3), .reg_partial_sum(spare_reg_psum_25_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_4( .activation_in(spare_reg_activation_25_3), .weight_in(spare_reg_weight_24_4), .partial_sum_in(spare_reg_psum_24_4), .reg_activation(spare_reg_activation_25_4), .reg_weight(spare_reg_weight_25_4), .reg_partial_sum(spare_reg_psum_25_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_5( .activation_in(spare_reg_activation_25_4), .weight_in(spare_reg_weight_24_5), .partial_sum_in(spare_reg_psum_24_5), .reg_activation(spare_reg_activation_25_5), .reg_weight(spare_reg_weight_25_5), .reg_partial_sum(spare_reg_psum_25_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_6( .activation_in(spare_reg_activation_25_5), .weight_in(spare_reg_weight_24_6), .partial_sum_in(spare_reg_psum_24_6), .reg_activation(spare_reg_activation_25_6), .reg_weight(spare_reg_weight_25_6), .reg_partial_sum(spare_reg_psum_25_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_7( .activation_in(spare_reg_activation_25_6), .weight_in(spare_reg_weight_24_7), .partial_sum_in(spare_reg_psum_24_7), .reg_activation(spare_reg_activation_25_7), .reg_weight(spare_reg_weight_25_7), .reg_partial_sum(spare_reg_psum_25_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_8( .activation_in(spare_reg_activation_25_7), .weight_in(spare_reg_weight_24_8), .partial_sum_in(spare_reg_psum_24_8), .reg_activation(spare_reg_activation_25_8), .reg_weight(spare_reg_weight_25_8), .reg_partial_sum(spare_reg_psum_25_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_9( .activation_in(spare_reg_activation_25_8), .weight_in(spare_reg_weight_24_9), .partial_sum_in(spare_reg_psum_24_9), .reg_activation(spare_reg_activation_25_9), .reg_weight(spare_reg_weight_25_9), .reg_partial_sum(spare_reg_psum_25_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_10( .activation_in(spare_reg_activation_25_9), .weight_in(spare_reg_weight_24_10), .partial_sum_in(spare_reg_psum_24_10), .reg_activation(spare_reg_activation_25_10), .reg_weight(spare_reg_weight_25_10), .reg_partial_sum(spare_reg_psum_25_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_11( .activation_in(spare_reg_activation_25_10), .weight_in(spare_reg_weight_24_11), .partial_sum_in(spare_reg_psum_24_11), .reg_activation(spare_reg_activation_25_11), .reg_weight(spare_reg_weight_25_11), .reg_partial_sum(spare_reg_psum_25_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_12( .activation_in(spare_reg_activation_25_11), .weight_in(spare_reg_weight_24_12), .partial_sum_in(spare_reg_psum_24_12), .reg_activation(spare_reg_activation_25_12), .reg_weight(spare_reg_weight_25_12), .reg_partial_sum(spare_reg_psum_25_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_13( .activation_in(spare_reg_activation_25_12), .weight_in(spare_reg_weight_24_13), .partial_sum_in(spare_reg_psum_24_13), .reg_activation(spare_reg_activation_25_13), .reg_weight(spare_reg_weight_25_13), .reg_partial_sum(spare_reg_psum_25_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_14( .activation_in(spare_reg_activation_25_13), .weight_in(spare_reg_weight_24_14), .partial_sum_in(spare_reg_psum_24_14), .reg_activation(spare_reg_activation_25_14), .reg_weight(spare_reg_weight_25_14), .reg_partial_sum(spare_reg_psum_25_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_15( .activation_in(spare_reg_activation_25_14), .weight_in(spare_reg_weight_24_15), .partial_sum_in(spare_reg_psum_24_15), .reg_activation(spare_reg_activation_25_15), .reg_weight(spare_reg_weight_25_15), .reg_partial_sum(spare_reg_psum_25_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_16( .activation_in(spare_reg_activation_25_15), .weight_in(spare_reg_weight_24_16), .partial_sum_in(spare_reg_psum_24_16), .reg_activation(spare_reg_activation_25_16), .reg_weight(spare_reg_weight_25_16), .reg_partial_sum(spare_reg_psum_25_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_17( .activation_in(spare_reg_activation_25_16), .weight_in(spare_reg_weight_24_17), .partial_sum_in(spare_reg_psum_24_17), .reg_activation(spare_reg_activation_25_17), .reg_weight(spare_reg_weight_25_17), .reg_partial_sum(spare_reg_psum_25_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_18( .activation_in(spare_reg_activation_25_17), .weight_in(spare_reg_weight_24_18), .partial_sum_in(spare_reg_psum_24_18), .reg_activation(spare_reg_activation_25_18), .reg_weight(spare_reg_weight_25_18), .reg_partial_sum(spare_reg_psum_25_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_19( .activation_in(spare_reg_activation_25_18), .weight_in(spare_reg_weight_24_19), .partial_sum_in(spare_reg_psum_24_19), .reg_activation(spare_reg_activation_25_19), .reg_weight(spare_reg_weight_25_19), .reg_partial_sum(spare_reg_psum_25_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_20( .activation_in(spare_reg_activation_25_19), .weight_in(spare_reg_weight_24_20), .partial_sum_in(spare_reg_psum_24_20), .reg_activation(spare_reg_activation_25_20), .reg_weight(spare_reg_weight_25_20), .reg_partial_sum(spare_reg_psum_25_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_21( .activation_in(spare_reg_activation_25_20), .weight_in(spare_reg_weight_24_21), .partial_sum_in(spare_reg_psum_24_21), .reg_activation(spare_reg_activation_25_21), .reg_weight(spare_reg_weight_25_21), .reg_partial_sum(spare_reg_psum_25_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_22( .activation_in(spare_reg_activation_25_21), .weight_in(spare_reg_weight_24_22), .partial_sum_in(spare_reg_psum_24_22), .reg_activation(spare_reg_activation_25_22), .reg_weight(spare_reg_weight_25_22), .reg_partial_sum(spare_reg_psum_25_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_23( .activation_in(spare_reg_activation_25_22), .weight_in(spare_reg_weight_24_23), .partial_sum_in(spare_reg_psum_24_23), .reg_activation(spare_reg_activation_25_23), .reg_weight(spare_reg_weight_25_23), .reg_partial_sum(spare_reg_psum_25_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_24( .activation_in(spare_reg_activation_25_23), .weight_in(spare_reg_weight_24_24), .partial_sum_in(spare_reg_psum_24_24), .reg_activation(spare_reg_activation_25_24), .reg_weight(spare_reg_weight_25_24), .reg_partial_sum(spare_reg_psum_25_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_25( .activation_in(spare_reg_activation_25_24), .weight_in(spare_reg_weight_24_25), .partial_sum_in(spare_reg_psum_24_25), .reg_activation(spare_reg_activation_25_25), .reg_weight(spare_reg_weight_25_25), .reg_partial_sum(spare_reg_psum_25_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_26( .activation_in(spare_reg_activation_25_25), .weight_in(spare_reg_weight_24_26), .partial_sum_in(spare_reg_psum_24_26), .reg_activation(spare_reg_activation_25_26), .reg_weight(spare_reg_weight_25_26), .reg_partial_sum(spare_reg_psum_25_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_27( .activation_in(spare_reg_activation_25_26), .weight_in(spare_reg_weight_24_27), .partial_sum_in(spare_reg_psum_24_27), .reg_activation(spare_reg_activation_25_27), .reg_weight(spare_reg_weight_25_27), .reg_partial_sum(spare_reg_psum_25_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_28( .activation_in(spare_reg_activation_25_27), .weight_in(spare_reg_weight_24_28), .partial_sum_in(spare_reg_psum_24_28), .reg_activation(spare_reg_activation_25_28), .reg_weight(spare_reg_weight_25_28), .reg_partial_sum(spare_reg_psum_25_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_29( .activation_in(spare_reg_activation_25_28), .weight_in(spare_reg_weight_24_29), .partial_sum_in(spare_reg_psum_24_29), .reg_activation(spare_reg_activation_25_29), .reg_weight(spare_reg_weight_25_29), .reg_partial_sum(spare_reg_psum_25_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_30( .activation_in(spare_reg_activation_25_29), .weight_in(spare_reg_weight_24_30), .partial_sum_in(spare_reg_psum_24_30), .reg_activation(spare_reg_activation_25_30), .reg_weight(spare_reg_weight_25_30), .reg_partial_sum(spare_reg_psum_25_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X25_31( .activation_in(spare_reg_activation_25_30), .weight_in(spare_reg_weight_24_31), .partial_sum_in(spare_reg_psum_24_31), .reg_weight(spare_reg_weight_25_31), .reg_partial_sum(spare_reg_psum_25_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_0( .activation_in(in_activation_26), .weight_in(spare_reg_weight_25_0), .partial_sum_in(spare_reg_psum_25_0), .reg_activation(spare_reg_activation_26_0), .reg_weight(spare_reg_weight_26_0), .reg_partial_sum(spare_reg_psum_26_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_1( .activation_in(spare_reg_activation_26_0), .weight_in(spare_reg_weight_25_1), .partial_sum_in(spare_reg_psum_25_1), .reg_activation(spare_reg_activation_26_1), .reg_weight(spare_reg_weight_26_1), .reg_partial_sum(spare_reg_psum_26_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_2( .activation_in(spare_reg_activation_26_1), .weight_in(spare_reg_weight_25_2), .partial_sum_in(spare_reg_psum_25_2), .reg_activation(spare_reg_activation_26_2), .reg_weight(spare_reg_weight_26_2), .reg_partial_sum(spare_reg_psum_26_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_3( .activation_in(spare_reg_activation_26_2), .weight_in(spare_reg_weight_25_3), .partial_sum_in(spare_reg_psum_25_3), .reg_activation(spare_reg_activation_26_3), .reg_weight(spare_reg_weight_26_3), .reg_partial_sum(spare_reg_psum_26_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_4( .activation_in(spare_reg_activation_26_3), .weight_in(spare_reg_weight_25_4), .partial_sum_in(spare_reg_psum_25_4), .reg_activation(spare_reg_activation_26_4), .reg_weight(spare_reg_weight_26_4), .reg_partial_sum(spare_reg_psum_26_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_5( .activation_in(spare_reg_activation_26_4), .weight_in(spare_reg_weight_25_5), .partial_sum_in(spare_reg_psum_25_5), .reg_activation(spare_reg_activation_26_5), .reg_weight(spare_reg_weight_26_5), .reg_partial_sum(spare_reg_psum_26_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_6( .activation_in(spare_reg_activation_26_5), .weight_in(spare_reg_weight_25_6), .partial_sum_in(spare_reg_psum_25_6), .reg_activation(spare_reg_activation_26_6), .reg_weight(spare_reg_weight_26_6), .reg_partial_sum(spare_reg_psum_26_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_7( .activation_in(spare_reg_activation_26_6), .weight_in(spare_reg_weight_25_7), .partial_sum_in(spare_reg_psum_25_7), .reg_activation(spare_reg_activation_26_7), .reg_weight(spare_reg_weight_26_7), .reg_partial_sum(spare_reg_psum_26_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_8( .activation_in(spare_reg_activation_26_7), .weight_in(spare_reg_weight_25_8), .partial_sum_in(spare_reg_psum_25_8), .reg_activation(spare_reg_activation_26_8), .reg_weight(spare_reg_weight_26_8), .reg_partial_sum(spare_reg_psum_26_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_9( .activation_in(spare_reg_activation_26_8), .weight_in(spare_reg_weight_25_9), .partial_sum_in(spare_reg_psum_25_9), .reg_activation(spare_reg_activation_26_9), .reg_weight(spare_reg_weight_26_9), .reg_partial_sum(spare_reg_psum_26_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_10( .activation_in(spare_reg_activation_26_9), .weight_in(spare_reg_weight_25_10), .partial_sum_in(spare_reg_psum_25_10), .reg_activation(spare_reg_activation_26_10), .reg_weight(spare_reg_weight_26_10), .reg_partial_sum(spare_reg_psum_26_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_11( .activation_in(spare_reg_activation_26_10), .weight_in(spare_reg_weight_25_11), .partial_sum_in(spare_reg_psum_25_11), .reg_activation(spare_reg_activation_26_11), .reg_weight(spare_reg_weight_26_11), .reg_partial_sum(spare_reg_psum_26_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_12( .activation_in(spare_reg_activation_26_11), .weight_in(spare_reg_weight_25_12), .partial_sum_in(spare_reg_psum_25_12), .reg_activation(spare_reg_activation_26_12), .reg_weight(spare_reg_weight_26_12), .reg_partial_sum(spare_reg_psum_26_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_13( .activation_in(spare_reg_activation_26_12), .weight_in(spare_reg_weight_25_13), .partial_sum_in(spare_reg_psum_25_13), .reg_activation(spare_reg_activation_26_13), .reg_weight(spare_reg_weight_26_13), .reg_partial_sum(spare_reg_psum_26_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_14( .activation_in(spare_reg_activation_26_13), .weight_in(spare_reg_weight_25_14), .partial_sum_in(spare_reg_psum_25_14), .reg_activation(spare_reg_activation_26_14), .reg_weight(spare_reg_weight_26_14), .reg_partial_sum(spare_reg_psum_26_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_15( .activation_in(spare_reg_activation_26_14), .weight_in(spare_reg_weight_25_15), .partial_sum_in(spare_reg_psum_25_15), .reg_activation(spare_reg_activation_26_15), .reg_weight(spare_reg_weight_26_15), .reg_partial_sum(spare_reg_psum_26_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_16( .activation_in(spare_reg_activation_26_15), .weight_in(spare_reg_weight_25_16), .partial_sum_in(spare_reg_psum_25_16), .reg_activation(spare_reg_activation_26_16), .reg_weight(spare_reg_weight_26_16), .reg_partial_sum(spare_reg_psum_26_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_17( .activation_in(spare_reg_activation_26_16), .weight_in(spare_reg_weight_25_17), .partial_sum_in(spare_reg_psum_25_17), .reg_activation(spare_reg_activation_26_17), .reg_weight(spare_reg_weight_26_17), .reg_partial_sum(spare_reg_psum_26_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_18( .activation_in(spare_reg_activation_26_17), .weight_in(spare_reg_weight_25_18), .partial_sum_in(spare_reg_psum_25_18), .reg_activation(spare_reg_activation_26_18), .reg_weight(spare_reg_weight_26_18), .reg_partial_sum(spare_reg_psum_26_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_19( .activation_in(spare_reg_activation_26_18), .weight_in(spare_reg_weight_25_19), .partial_sum_in(spare_reg_psum_25_19), .reg_activation(spare_reg_activation_26_19), .reg_weight(spare_reg_weight_26_19), .reg_partial_sum(spare_reg_psum_26_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_20( .activation_in(spare_reg_activation_26_19), .weight_in(spare_reg_weight_25_20), .partial_sum_in(spare_reg_psum_25_20), .reg_activation(spare_reg_activation_26_20), .reg_weight(spare_reg_weight_26_20), .reg_partial_sum(spare_reg_psum_26_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_21( .activation_in(spare_reg_activation_26_20), .weight_in(spare_reg_weight_25_21), .partial_sum_in(spare_reg_psum_25_21), .reg_activation(spare_reg_activation_26_21), .reg_weight(spare_reg_weight_26_21), .reg_partial_sum(spare_reg_psum_26_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_22( .activation_in(spare_reg_activation_26_21), .weight_in(spare_reg_weight_25_22), .partial_sum_in(spare_reg_psum_25_22), .reg_activation(spare_reg_activation_26_22), .reg_weight(spare_reg_weight_26_22), .reg_partial_sum(spare_reg_psum_26_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_23( .activation_in(spare_reg_activation_26_22), .weight_in(spare_reg_weight_25_23), .partial_sum_in(spare_reg_psum_25_23), .reg_activation(spare_reg_activation_26_23), .reg_weight(spare_reg_weight_26_23), .reg_partial_sum(spare_reg_psum_26_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_24( .activation_in(spare_reg_activation_26_23), .weight_in(spare_reg_weight_25_24), .partial_sum_in(spare_reg_psum_25_24), .reg_activation(spare_reg_activation_26_24), .reg_weight(spare_reg_weight_26_24), .reg_partial_sum(spare_reg_psum_26_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_25( .activation_in(spare_reg_activation_26_24), .weight_in(spare_reg_weight_25_25), .partial_sum_in(spare_reg_psum_25_25), .reg_activation(spare_reg_activation_26_25), .reg_weight(spare_reg_weight_26_25), .reg_partial_sum(spare_reg_psum_26_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_26( .activation_in(spare_reg_activation_26_25), .weight_in(spare_reg_weight_25_26), .partial_sum_in(spare_reg_psum_25_26), .reg_activation(spare_reg_activation_26_26), .reg_weight(spare_reg_weight_26_26), .reg_partial_sum(spare_reg_psum_26_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_27( .activation_in(spare_reg_activation_26_26), .weight_in(spare_reg_weight_25_27), .partial_sum_in(spare_reg_psum_25_27), .reg_activation(spare_reg_activation_26_27), .reg_weight(spare_reg_weight_26_27), .reg_partial_sum(spare_reg_psum_26_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_28( .activation_in(spare_reg_activation_26_27), .weight_in(spare_reg_weight_25_28), .partial_sum_in(spare_reg_psum_25_28), .reg_activation(spare_reg_activation_26_28), .reg_weight(spare_reg_weight_26_28), .reg_partial_sum(spare_reg_psum_26_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_29( .activation_in(spare_reg_activation_26_28), .weight_in(spare_reg_weight_25_29), .partial_sum_in(spare_reg_psum_25_29), .reg_activation(spare_reg_activation_26_29), .reg_weight(spare_reg_weight_26_29), .reg_partial_sum(spare_reg_psum_26_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_30( .activation_in(spare_reg_activation_26_29), .weight_in(spare_reg_weight_25_30), .partial_sum_in(spare_reg_psum_25_30), .reg_activation(spare_reg_activation_26_30), .reg_weight(spare_reg_weight_26_30), .reg_partial_sum(spare_reg_psum_26_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X26_31( .activation_in(spare_reg_activation_26_30), .weight_in(spare_reg_weight_25_31), .partial_sum_in(spare_reg_psum_25_31), .reg_weight(spare_reg_weight_26_31), .reg_partial_sum(spare_reg_psum_26_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_0( .activation_in(in_activation_27), .weight_in(spare_reg_weight_26_0), .partial_sum_in(spare_reg_psum_26_0), .reg_activation(spare_reg_activation_27_0), .reg_weight(spare_reg_weight_27_0), .reg_partial_sum(spare_reg_psum_27_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_1( .activation_in(spare_reg_activation_27_0), .weight_in(spare_reg_weight_26_1), .partial_sum_in(spare_reg_psum_26_1), .reg_activation(spare_reg_activation_27_1), .reg_weight(spare_reg_weight_27_1), .reg_partial_sum(spare_reg_psum_27_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_2( .activation_in(spare_reg_activation_27_1), .weight_in(spare_reg_weight_26_2), .partial_sum_in(spare_reg_psum_26_2), .reg_activation(spare_reg_activation_27_2), .reg_weight(spare_reg_weight_27_2), .reg_partial_sum(spare_reg_psum_27_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_3( .activation_in(spare_reg_activation_27_2), .weight_in(spare_reg_weight_26_3), .partial_sum_in(spare_reg_psum_26_3), .reg_activation(spare_reg_activation_27_3), .reg_weight(spare_reg_weight_27_3), .reg_partial_sum(spare_reg_psum_27_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_4( .activation_in(spare_reg_activation_27_3), .weight_in(spare_reg_weight_26_4), .partial_sum_in(spare_reg_psum_26_4), .reg_activation(spare_reg_activation_27_4), .reg_weight(spare_reg_weight_27_4), .reg_partial_sum(spare_reg_psum_27_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_5( .activation_in(spare_reg_activation_27_4), .weight_in(spare_reg_weight_26_5), .partial_sum_in(spare_reg_psum_26_5), .reg_activation(spare_reg_activation_27_5), .reg_weight(spare_reg_weight_27_5), .reg_partial_sum(spare_reg_psum_27_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_6( .activation_in(spare_reg_activation_27_5), .weight_in(spare_reg_weight_26_6), .partial_sum_in(spare_reg_psum_26_6), .reg_activation(spare_reg_activation_27_6), .reg_weight(spare_reg_weight_27_6), .reg_partial_sum(spare_reg_psum_27_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_7( .activation_in(spare_reg_activation_27_6), .weight_in(spare_reg_weight_26_7), .partial_sum_in(spare_reg_psum_26_7), .reg_activation(spare_reg_activation_27_7), .reg_weight(spare_reg_weight_27_7), .reg_partial_sum(spare_reg_psum_27_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_8( .activation_in(spare_reg_activation_27_7), .weight_in(spare_reg_weight_26_8), .partial_sum_in(spare_reg_psum_26_8), .reg_activation(spare_reg_activation_27_8), .reg_weight(spare_reg_weight_27_8), .reg_partial_sum(spare_reg_psum_27_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_9( .activation_in(spare_reg_activation_27_8), .weight_in(spare_reg_weight_26_9), .partial_sum_in(spare_reg_psum_26_9), .reg_activation(spare_reg_activation_27_9), .reg_weight(spare_reg_weight_27_9), .reg_partial_sum(spare_reg_psum_27_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_10( .activation_in(spare_reg_activation_27_9), .weight_in(spare_reg_weight_26_10), .partial_sum_in(spare_reg_psum_26_10), .reg_activation(spare_reg_activation_27_10), .reg_weight(spare_reg_weight_27_10), .reg_partial_sum(spare_reg_psum_27_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_11( .activation_in(spare_reg_activation_27_10), .weight_in(spare_reg_weight_26_11), .partial_sum_in(spare_reg_psum_26_11), .reg_activation(spare_reg_activation_27_11), .reg_weight(spare_reg_weight_27_11), .reg_partial_sum(spare_reg_psum_27_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_12( .activation_in(spare_reg_activation_27_11), .weight_in(spare_reg_weight_26_12), .partial_sum_in(spare_reg_psum_26_12), .reg_activation(spare_reg_activation_27_12), .reg_weight(spare_reg_weight_27_12), .reg_partial_sum(spare_reg_psum_27_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_13( .activation_in(spare_reg_activation_27_12), .weight_in(spare_reg_weight_26_13), .partial_sum_in(spare_reg_psum_26_13), .reg_activation(spare_reg_activation_27_13), .reg_weight(spare_reg_weight_27_13), .reg_partial_sum(spare_reg_psum_27_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_14( .activation_in(spare_reg_activation_27_13), .weight_in(spare_reg_weight_26_14), .partial_sum_in(spare_reg_psum_26_14), .reg_activation(spare_reg_activation_27_14), .reg_weight(spare_reg_weight_27_14), .reg_partial_sum(spare_reg_psum_27_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_15( .activation_in(spare_reg_activation_27_14), .weight_in(spare_reg_weight_26_15), .partial_sum_in(spare_reg_psum_26_15), .reg_activation(spare_reg_activation_27_15), .reg_weight(spare_reg_weight_27_15), .reg_partial_sum(spare_reg_psum_27_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_16( .activation_in(spare_reg_activation_27_15), .weight_in(spare_reg_weight_26_16), .partial_sum_in(spare_reg_psum_26_16), .reg_activation(spare_reg_activation_27_16), .reg_weight(spare_reg_weight_27_16), .reg_partial_sum(spare_reg_psum_27_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_17( .activation_in(spare_reg_activation_27_16), .weight_in(spare_reg_weight_26_17), .partial_sum_in(spare_reg_psum_26_17), .reg_activation(spare_reg_activation_27_17), .reg_weight(spare_reg_weight_27_17), .reg_partial_sum(spare_reg_psum_27_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_18( .activation_in(spare_reg_activation_27_17), .weight_in(spare_reg_weight_26_18), .partial_sum_in(spare_reg_psum_26_18), .reg_activation(spare_reg_activation_27_18), .reg_weight(spare_reg_weight_27_18), .reg_partial_sum(spare_reg_psum_27_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_19( .activation_in(spare_reg_activation_27_18), .weight_in(spare_reg_weight_26_19), .partial_sum_in(spare_reg_psum_26_19), .reg_activation(spare_reg_activation_27_19), .reg_weight(spare_reg_weight_27_19), .reg_partial_sum(spare_reg_psum_27_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_20( .activation_in(spare_reg_activation_27_19), .weight_in(spare_reg_weight_26_20), .partial_sum_in(spare_reg_psum_26_20), .reg_activation(spare_reg_activation_27_20), .reg_weight(spare_reg_weight_27_20), .reg_partial_sum(spare_reg_psum_27_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_21( .activation_in(spare_reg_activation_27_20), .weight_in(spare_reg_weight_26_21), .partial_sum_in(spare_reg_psum_26_21), .reg_activation(spare_reg_activation_27_21), .reg_weight(spare_reg_weight_27_21), .reg_partial_sum(spare_reg_psum_27_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_22( .activation_in(spare_reg_activation_27_21), .weight_in(spare_reg_weight_26_22), .partial_sum_in(spare_reg_psum_26_22), .reg_activation(spare_reg_activation_27_22), .reg_weight(spare_reg_weight_27_22), .reg_partial_sum(spare_reg_psum_27_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_23( .activation_in(spare_reg_activation_27_22), .weight_in(spare_reg_weight_26_23), .partial_sum_in(spare_reg_psum_26_23), .reg_activation(spare_reg_activation_27_23), .reg_weight(spare_reg_weight_27_23), .reg_partial_sum(spare_reg_psum_27_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_24( .activation_in(spare_reg_activation_27_23), .weight_in(spare_reg_weight_26_24), .partial_sum_in(spare_reg_psum_26_24), .reg_activation(spare_reg_activation_27_24), .reg_weight(spare_reg_weight_27_24), .reg_partial_sum(spare_reg_psum_27_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_25( .activation_in(spare_reg_activation_27_24), .weight_in(spare_reg_weight_26_25), .partial_sum_in(spare_reg_psum_26_25), .reg_activation(spare_reg_activation_27_25), .reg_weight(spare_reg_weight_27_25), .reg_partial_sum(spare_reg_psum_27_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_26( .activation_in(spare_reg_activation_27_25), .weight_in(spare_reg_weight_26_26), .partial_sum_in(spare_reg_psum_26_26), .reg_activation(spare_reg_activation_27_26), .reg_weight(spare_reg_weight_27_26), .reg_partial_sum(spare_reg_psum_27_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_27( .activation_in(spare_reg_activation_27_26), .weight_in(spare_reg_weight_26_27), .partial_sum_in(spare_reg_psum_26_27), .reg_activation(spare_reg_activation_27_27), .reg_weight(spare_reg_weight_27_27), .reg_partial_sum(spare_reg_psum_27_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_28( .activation_in(spare_reg_activation_27_27), .weight_in(spare_reg_weight_26_28), .partial_sum_in(spare_reg_psum_26_28), .reg_activation(spare_reg_activation_27_28), .reg_weight(spare_reg_weight_27_28), .reg_partial_sum(spare_reg_psum_27_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_29( .activation_in(spare_reg_activation_27_28), .weight_in(spare_reg_weight_26_29), .partial_sum_in(spare_reg_psum_26_29), .reg_activation(spare_reg_activation_27_29), .reg_weight(spare_reg_weight_27_29), .reg_partial_sum(spare_reg_psum_27_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_30( .activation_in(spare_reg_activation_27_29), .weight_in(spare_reg_weight_26_30), .partial_sum_in(spare_reg_psum_26_30), .reg_activation(spare_reg_activation_27_30), .reg_weight(spare_reg_weight_27_30), .reg_partial_sum(spare_reg_psum_27_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X27_31( .activation_in(spare_reg_activation_27_30), .weight_in(spare_reg_weight_26_31), .partial_sum_in(spare_reg_psum_26_31), .reg_weight(spare_reg_weight_27_31), .reg_partial_sum(spare_reg_psum_27_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_0( .activation_in(in_activation_28), .weight_in(spare_reg_weight_27_0), .partial_sum_in(spare_reg_psum_27_0), .reg_activation(spare_reg_activation_28_0), .reg_weight(spare_reg_weight_28_0), .reg_partial_sum(spare_reg_psum_28_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_1( .activation_in(spare_reg_activation_28_0), .weight_in(spare_reg_weight_27_1), .partial_sum_in(spare_reg_psum_27_1), .reg_activation(spare_reg_activation_28_1), .reg_weight(spare_reg_weight_28_1), .reg_partial_sum(spare_reg_psum_28_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_2( .activation_in(spare_reg_activation_28_1), .weight_in(spare_reg_weight_27_2), .partial_sum_in(spare_reg_psum_27_2), .reg_activation(spare_reg_activation_28_2), .reg_weight(spare_reg_weight_28_2), .reg_partial_sum(spare_reg_psum_28_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_3( .activation_in(spare_reg_activation_28_2), .weight_in(spare_reg_weight_27_3), .partial_sum_in(spare_reg_psum_27_3), .reg_activation(spare_reg_activation_28_3), .reg_weight(spare_reg_weight_28_3), .reg_partial_sum(spare_reg_psum_28_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_4( .activation_in(spare_reg_activation_28_3), .weight_in(spare_reg_weight_27_4), .partial_sum_in(spare_reg_psum_27_4), .reg_activation(spare_reg_activation_28_4), .reg_weight(spare_reg_weight_28_4), .reg_partial_sum(spare_reg_psum_28_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_5( .activation_in(spare_reg_activation_28_4), .weight_in(spare_reg_weight_27_5), .partial_sum_in(spare_reg_psum_27_5), .reg_activation(spare_reg_activation_28_5), .reg_weight(spare_reg_weight_28_5), .reg_partial_sum(spare_reg_psum_28_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_6( .activation_in(spare_reg_activation_28_5), .weight_in(spare_reg_weight_27_6), .partial_sum_in(spare_reg_psum_27_6), .reg_activation(spare_reg_activation_28_6), .reg_weight(spare_reg_weight_28_6), .reg_partial_sum(spare_reg_psum_28_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_7( .activation_in(spare_reg_activation_28_6), .weight_in(spare_reg_weight_27_7), .partial_sum_in(spare_reg_psum_27_7), .reg_activation(spare_reg_activation_28_7), .reg_weight(spare_reg_weight_28_7), .reg_partial_sum(spare_reg_psum_28_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_8( .activation_in(spare_reg_activation_28_7), .weight_in(spare_reg_weight_27_8), .partial_sum_in(spare_reg_psum_27_8), .reg_activation(spare_reg_activation_28_8), .reg_weight(spare_reg_weight_28_8), .reg_partial_sum(spare_reg_psum_28_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_9( .activation_in(spare_reg_activation_28_8), .weight_in(spare_reg_weight_27_9), .partial_sum_in(spare_reg_psum_27_9), .reg_activation(spare_reg_activation_28_9), .reg_weight(spare_reg_weight_28_9), .reg_partial_sum(spare_reg_psum_28_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_10( .activation_in(spare_reg_activation_28_9), .weight_in(spare_reg_weight_27_10), .partial_sum_in(spare_reg_psum_27_10), .reg_activation(spare_reg_activation_28_10), .reg_weight(spare_reg_weight_28_10), .reg_partial_sum(spare_reg_psum_28_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_11( .activation_in(spare_reg_activation_28_10), .weight_in(spare_reg_weight_27_11), .partial_sum_in(spare_reg_psum_27_11), .reg_activation(spare_reg_activation_28_11), .reg_weight(spare_reg_weight_28_11), .reg_partial_sum(spare_reg_psum_28_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_12( .activation_in(spare_reg_activation_28_11), .weight_in(spare_reg_weight_27_12), .partial_sum_in(spare_reg_psum_27_12), .reg_activation(spare_reg_activation_28_12), .reg_weight(spare_reg_weight_28_12), .reg_partial_sum(spare_reg_psum_28_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_13( .activation_in(spare_reg_activation_28_12), .weight_in(spare_reg_weight_27_13), .partial_sum_in(spare_reg_psum_27_13), .reg_activation(spare_reg_activation_28_13), .reg_weight(spare_reg_weight_28_13), .reg_partial_sum(spare_reg_psum_28_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_14( .activation_in(spare_reg_activation_28_13), .weight_in(spare_reg_weight_27_14), .partial_sum_in(spare_reg_psum_27_14), .reg_activation(spare_reg_activation_28_14), .reg_weight(spare_reg_weight_28_14), .reg_partial_sum(spare_reg_psum_28_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_15( .activation_in(spare_reg_activation_28_14), .weight_in(spare_reg_weight_27_15), .partial_sum_in(spare_reg_psum_27_15), .reg_activation(spare_reg_activation_28_15), .reg_weight(spare_reg_weight_28_15), .reg_partial_sum(spare_reg_psum_28_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_16( .activation_in(spare_reg_activation_28_15), .weight_in(spare_reg_weight_27_16), .partial_sum_in(spare_reg_psum_27_16), .reg_activation(spare_reg_activation_28_16), .reg_weight(spare_reg_weight_28_16), .reg_partial_sum(spare_reg_psum_28_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_17( .activation_in(spare_reg_activation_28_16), .weight_in(spare_reg_weight_27_17), .partial_sum_in(spare_reg_psum_27_17), .reg_activation(spare_reg_activation_28_17), .reg_weight(spare_reg_weight_28_17), .reg_partial_sum(spare_reg_psum_28_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_18( .activation_in(spare_reg_activation_28_17), .weight_in(spare_reg_weight_27_18), .partial_sum_in(spare_reg_psum_27_18), .reg_activation(spare_reg_activation_28_18), .reg_weight(spare_reg_weight_28_18), .reg_partial_sum(spare_reg_psum_28_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_19( .activation_in(spare_reg_activation_28_18), .weight_in(spare_reg_weight_27_19), .partial_sum_in(spare_reg_psum_27_19), .reg_activation(spare_reg_activation_28_19), .reg_weight(spare_reg_weight_28_19), .reg_partial_sum(spare_reg_psum_28_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_20( .activation_in(spare_reg_activation_28_19), .weight_in(spare_reg_weight_27_20), .partial_sum_in(spare_reg_psum_27_20), .reg_activation(spare_reg_activation_28_20), .reg_weight(spare_reg_weight_28_20), .reg_partial_sum(spare_reg_psum_28_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_21( .activation_in(spare_reg_activation_28_20), .weight_in(spare_reg_weight_27_21), .partial_sum_in(spare_reg_psum_27_21), .reg_activation(spare_reg_activation_28_21), .reg_weight(spare_reg_weight_28_21), .reg_partial_sum(spare_reg_psum_28_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_22( .activation_in(spare_reg_activation_28_21), .weight_in(spare_reg_weight_27_22), .partial_sum_in(spare_reg_psum_27_22), .reg_activation(spare_reg_activation_28_22), .reg_weight(spare_reg_weight_28_22), .reg_partial_sum(spare_reg_psum_28_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_23( .activation_in(spare_reg_activation_28_22), .weight_in(spare_reg_weight_27_23), .partial_sum_in(spare_reg_psum_27_23), .reg_activation(spare_reg_activation_28_23), .reg_weight(spare_reg_weight_28_23), .reg_partial_sum(spare_reg_psum_28_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_24( .activation_in(spare_reg_activation_28_23), .weight_in(spare_reg_weight_27_24), .partial_sum_in(spare_reg_psum_27_24), .reg_activation(spare_reg_activation_28_24), .reg_weight(spare_reg_weight_28_24), .reg_partial_sum(spare_reg_psum_28_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_25( .activation_in(spare_reg_activation_28_24), .weight_in(spare_reg_weight_27_25), .partial_sum_in(spare_reg_psum_27_25), .reg_activation(spare_reg_activation_28_25), .reg_weight(spare_reg_weight_28_25), .reg_partial_sum(spare_reg_psum_28_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_26( .activation_in(spare_reg_activation_28_25), .weight_in(spare_reg_weight_27_26), .partial_sum_in(spare_reg_psum_27_26), .reg_activation(spare_reg_activation_28_26), .reg_weight(spare_reg_weight_28_26), .reg_partial_sum(spare_reg_psum_28_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_27( .activation_in(spare_reg_activation_28_26), .weight_in(spare_reg_weight_27_27), .partial_sum_in(spare_reg_psum_27_27), .reg_activation(spare_reg_activation_28_27), .reg_weight(spare_reg_weight_28_27), .reg_partial_sum(spare_reg_psum_28_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_28( .activation_in(spare_reg_activation_28_27), .weight_in(spare_reg_weight_27_28), .partial_sum_in(spare_reg_psum_27_28), .reg_activation(spare_reg_activation_28_28), .reg_weight(spare_reg_weight_28_28), .reg_partial_sum(spare_reg_psum_28_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_29( .activation_in(spare_reg_activation_28_28), .weight_in(spare_reg_weight_27_29), .partial_sum_in(spare_reg_psum_27_29), .reg_activation(spare_reg_activation_28_29), .reg_weight(spare_reg_weight_28_29), .reg_partial_sum(spare_reg_psum_28_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_30( .activation_in(spare_reg_activation_28_29), .weight_in(spare_reg_weight_27_30), .partial_sum_in(spare_reg_psum_27_30), .reg_activation(spare_reg_activation_28_30), .reg_weight(spare_reg_weight_28_30), .reg_partial_sum(spare_reg_psum_28_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X28_31( .activation_in(spare_reg_activation_28_30), .weight_in(spare_reg_weight_27_31), .partial_sum_in(spare_reg_psum_27_31), .reg_weight(spare_reg_weight_28_31), .reg_partial_sum(spare_reg_psum_28_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_0( .activation_in(in_activation_29), .weight_in(spare_reg_weight_28_0), .partial_sum_in(spare_reg_psum_28_0), .reg_activation(spare_reg_activation_29_0), .reg_weight(spare_reg_weight_29_0), .reg_partial_sum(spare_reg_psum_29_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_1( .activation_in(spare_reg_activation_29_0), .weight_in(spare_reg_weight_28_1), .partial_sum_in(spare_reg_psum_28_1), .reg_activation(spare_reg_activation_29_1), .reg_weight(spare_reg_weight_29_1), .reg_partial_sum(spare_reg_psum_29_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_2( .activation_in(spare_reg_activation_29_1), .weight_in(spare_reg_weight_28_2), .partial_sum_in(spare_reg_psum_28_2), .reg_activation(spare_reg_activation_29_2), .reg_weight(spare_reg_weight_29_2), .reg_partial_sum(spare_reg_psum_29_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_3( .activation_in(spare_reg_activation_29_2), .weight_in(spare_reg_weight_28_3), .partial_sum_in(spare_reg_psum_28_3), .reg_activation(spare_reg_activation_29_3), .reg_weight(spare_reg_weight_29_3), .reg_partial_sum(spare_reg_psum_29_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_4( .activation_in(spare_reg_activation_29_3), .weight_in(spare_reg_weight_28_4), .partial_sum_in(spare_reg_psum_28_4), .reg_activation(spare_reg_activation_29_4), .reg_weight(spare_reg_weight_29_4), .reg_partial_sum(spare_reg_psum_29_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_5( .activation_in(spare_reg_activation_29_4), .weight_in(spare_reg_weight_28_5), .partial_sum_in(spare_reg_psum_28_5), .reg_activation(spare_reg_activation_29_5), .reg_weight(spare_reg_weight_29_5), .reg_partial_sum(spare_reg_psum_29_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_6( .activation_in(spare_reg_activation_29_5), .weight_in(spare_reg_weight_28_6), .partial_sum_in(spare_reg_psum_28_6), .reg_activation(spare_reg_activation_29_6), .reg_weight(spare_reg_weight_29_6), .reg_partial_sum(spare_reg_psum_29_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_7( .activation_in(spare_reg_activation_29_6), .weight_in(spare_reg_weight_28_7), .partial_sum_in(spare_reg_psum_28_7), .reg_activation(spare_reg_activation_29_7), .reg_weight(spare_reg_weight_29_7), .reg_partial_sum(spare_reg_psum_29_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_8( .activation_in(spare_reg_activation_29_7), .weight_in(spare_reg_weight_28_8), .partial_sum_in(spare_reg_psum_28_8), .reg_activation(spare_reg_activation_29_8), .reg_weight(spare_reg_weight_29_8), .reg_partial_sum(spare_reg_psum_29_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_9( .activation_in(spare_reg_activation_29_8), .weight_in(spare_reg_weight_28_9), .partial_sum_in(spare_reg_psum_28_9), .reg_activation(spare_reg_activation_29_9), .reg_weight(spare_reg_weight_29_9), .reg_partial_sum(spare_reg_psum_29_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_10( .activation_in(spare_reg_activation_29_9), .weight_in(spare_reg_weight_28_10), .partial_sum_in(spare_reg_psum_28_10), .reg_activation(spare_reg_activation_29_10), .reg_weight(spare_reg_weight_29_10), .reg_partial_sum(spare_reg_psum_29_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_11( .activation_in(spare_reg_activation_29_10), .weight_in(spare_reg_weight_28_11), .partial_sum_in(spare_reg_psum_28_11), .reg_activation(spare_reg_activation_29_11), .reg_weight(spare_reg_weight_29_11), .reg_partial_sum(spare_reg_psum_29_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_12( .activation_in(spare_reg_activation_29_11), .weight_in(spare_reg_weight_28_12), .partial_sum_in(spare_reg_psum_28_12), .reg_activation(spare_reg_activation_29_12), .reg_weight(spare_reg_weight_29_12), .reg_partial_sum(spare_reg_psum_29_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_13( .activation_in(spare_reg_activation_29_12), .weight_in(spare_reg_weight_28_13), .partial_sum_in(spare_reg_psum_28_13), .reg_activation(spare_reg_activation_29_13), .reg_weight(spare_reg_weight_29_13), .reg_partial_sum(spare_reg_psum_29_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_14( .activation_in(spare_reg_activation_29_13), .weight_in(spare_reg_weight_28_14), .partial_sum_in(spare_reg_psum_28_14), .reg_activation(spare_reg_activation_29_14), .reg_weight(spare_reg_weight_29_14), .reg_partial_sum(spare_reg_psum_29_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_15( .activation_in(spare_reg_activation_29_14), .weight_in(spare_reg_weight_28_15), .partial_sum_in(spare_reg_psum_28_15), .reg_activation(spare_reg_activation_29_15), .reg_weight(spare_reg_weight_29_15), .reg_partial_sum(spare_reg_psum_29_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_16( .activation_in(spare_reg_activation_29_15), .weight_in(spare_reg_weight_28_16), .partial_sum_in(spare_reg_psum_28_16), .reg_activation(spare_reg_activation_29_16), .reg_weight(spare_reg_weight_29_16), .reg_partial_sum(spare_reg_psum_29_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_17( .activation_in(spare_reg_activation_29_16), .weight_in(spare_reg_weight_28_17), .partial_sum_in(spare_reg_psum_28_17), .reg_activation(spare_reg_activation_29_17), .reg_weight(spare_reg_weight_29_17), .reg_partial_sum(spare_reg_psum_29_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_18( .activation_in(spare_reg_activation_29_17), .weight_in(spare_reg_weight_28_18), .partial_sum_in(spare_reg_psum_28_18), .reg_activation(spare_reg_activation_29_18), .reg_weight(spare_reg_weight_29_18), .reg_partial_sum(spare_reg_psum_29_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_19( .activation_in(spare_reg_activation_29_18), .weight_in(spare_reg_weight_28_19), .partial_sum_in(spare_reg_psum_28_19), .reg_activation(spare_reg_activation_29_19), .reg_weight(spare_reg_weight_29_19), .reg_partial_sum(spare_reg_psum_29_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_20( .activation_in(spare_reg_activation_29_19), .weight_in(spare_reg_weight_28_20), .partial_sum_in(spare_reg_psum_28_20), .reg_activation(spare_reg_activation_29_20), .reg_weight(spare_reg_weight_29_20), .reg_partial_sum(spare_reg_psum_29_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_21( .activation_in(spare_reg_activation_29_20), .weight_in(spare_reg_weight_28_21), .partial_sum_in(spare_reg_psum_28_21), .reg_activation(spare_reg_activation_29_21), .reg_weight(spare_reg_weight_29_21), .reg_partial_sum(spare_reg_psum_29_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_22( .activation_in(spare_reg_activation_29_21), .weight_in(spare_reg_weight_28_22), .partial_sum_in(spare_reg_psum_28_22), .reg_activation(spare_reg_activation_29_22), .reg_weight(spare_reg_weight_29_22), .reg_partial_sum(spare_reg_psum_29_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_23( .activation_in(spare_reg_activation_29_22), .weight_in(spare_reg_weight_28_23), .partial_sum_in(spare_reg_psum_28_23), .reg_activation(spare_reg_activation_29_23), .reg_weight(spare_reg_weight_29_23), .reg_partial_sum(spare_reg_psum_29_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_24( .activation_in(spare_reg_activation_29_23), .weight_in(spare_reg_weight_28_24), .partial_sum_in(spare_reg_psum_28_24), .reg_activation(spare_reg_activation_29_24), .reg_weight(spare_reg_weight_29_24), .reg_partial_sum(spare_reg_psum_29_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_25( .activation_in(spare_reg_activation_29_24), .weight_in(spare_reg_weight_28_25), .partial_sum_in(spare_reg_psum_28_25), .reg_activation(spare_reg_activation_29_25), .reg_weight(spare_reg_weight_29_25), .reg_partial_sum(spare_reg_psum_29_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_26( .activation_in(spare_reg_activation_29_25), .weight_in(spare_reg_weight_28_26), .partial_sum_in(spare_reg_psum_28_26), .reg_activation(spare_reg_activation_29_26), .reg_weight(spare_reg_weight_29_26), .reg_partial_sum(spare_reg_psum_29_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_27( .activation_in(spare_reg_activation_29_26), .weight_in(spare_reg_weight_28_27), .partial_sum_in(spare_reg_psum_28_27), .reg_activation(spare_reg_activation_29_27), .reg_weight(spare_reg_weight_29_27), .reg_partial_sum(spare_reg_psum_29_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_28( .activation_in(spare_reg_activation_29_27), .weight_in(spare_reg_weight_28_28), .partial_sum_in(spare_reg_psum_28_28), .reg_activation(spare_reg_activation_29_28), .reg_weight(spare_reg_weight_29_28), .reg_partial_sum(spare_reg_psum_29_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_29( .activation_in(spare_reg_activation_29_28), .weight_in(spare_reg_weight_28_29), .partial_sum_in(spare_reg_psum_28_29), .reg_activation(spare_reg_activation_29_29), .reg_weight(spare_reg_weight_29_29), .reg_partial_sum(spare_reg_psum_29_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_30( .activation_in(spare_reg_activation_29_29), .weight_in(spare_reg_weight_28_30), .partial_sum_in(spare_reg_psum_28_30), .reg_activation(spare_reg_activation_29_30), .reg_weight(spare_reg_weight_29_30), .reg_partial_sum(spare_reg_psum_29_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X29_31( .activation_in(spare_reg_activation_29_30), .weight_in(spare_reg_weight_28_31), .partial_sum_in(spare_reg_psum_28_31), .reg_weight(spare_reg_weight_29_31), .reg_partial_sum(spare_reg_psum_29_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_0( .activation_in(in_activation_30), .weight_in(spare_reg_weight_29_0), .partial_sum_in(spare_reg_psum_29_0), .reg_activation(spare_reg_activation_30_0), .reg_weight(spare_reg_weight_30_0), .reg_partial_sum(spare_reg_psum_30_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_1( .activation_in(spare_reg_activation_30_0), .weight_in(spare_reg_weight_29_1), .partial_sum_in(spare_reg_psum_29_1), .reg_activation(spare_reg_activation_30_1), .reg_weight(spare_reg_weight_30_1), .reg_partial_sum(spare_reg_psum_30_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_2( .activation_in(spare_reg_activation_30_1), .weight_in(spare_reg_weight_29_2), .partial_sum_in(spare_reg_psum_29_2), .reg_activation(spare_reg_activation_30_2), .reg_weight(spare_reg_weight_30_2), .reg_partial_sum(spare_reg_psum_30_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_3( .activation_in(spare_reg_activation_30_2), .weight_in(spare_reg_weight_29_3), .partial_sum_in(spare_reg_psum_29_3), .reg_activation(spare_reg_activation_30_3), .reg_weight(spare_reg_weight_30_3), .reg_partial_sum(spare_reg_psum_30_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_4( .activation_in(spare_reg_activation_30_3), .weight_in(spare_reg_weight_29_4), .partial_sum_in(spare_reg_psum_29_4), .reg_activation(spare_reg_activation_30_4), .reg_weight(spare_reg_weight_30_4), .reg_partial_sum(spare_reg_psum_30_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_5( .activation_in(spare_reg_activation_30_4), .weight_in(spare_reg_weight_29_5), .partial_sum_in(spare_reg_psum_29_5), .reg_activation(spare_reg_activation_30_5), .reg_weight(spare_reg_weight_30_5), .reg_partial_sum(spare_reg_psum_30_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_6( .activation_in(spare_reg_activation_30_5), .weight_in(spare_reg_weight_29_6), .partial_sum_in(spare_reg_psum_29_6), .reg_activation(spare_reg_activation_30_6), .reg_weight(spare_reg_weight_30_6), .reg_partial_sum(spare_reg_psum_30_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_7( .activation_in(spare_reg_activation_30_6), .weight_in(spare_reg_weight_29_7), .partial_sum_in(spare_reg_psum_29_7), .reg_activation(spare_reg_activation_30_7), .reg_weight(spare_reg_weight_30_7), .reg_partial_sum(spare_reg_psum_30_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_8( .activation_in(spare_reg_activation_30_7), .weight_in(spare_reg_weight_29_8), .partial_sum_in(spare_reg_psum_29_8), .reg_activation(spare_reg_activation_30_8), .reg_weight(spare_reg_weight_30_8), .reg_partial_sum(spare_reg_psum_30_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_9( .activation_in(spare_reg_activation_30_8), .weight_in(spare_reg_weight_29_9), .partial_sum_in(spare_reg_psum_29_9), .reg_activation(spare_reg_activation_30_9), .reg_weight(spare_reg_weight_30_9), .reg_partial_sum(spare_reg_psum_30_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_10( .activation_in(spare_reg_activation_30_9), .weight_in(spare_reg_weight_29_10), .partial_sum_in(spare_reg_psum_29_10), .reg_activation(spare_reg_activation_30_10), .reg_weight(spare_reg_weight_30_10), .reg_partial_sum(spare_reg_psum_30_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_11( .activation_in(spare_reg_activation_30_10), .weight_in(spare_reg_weight_29_11), .partial_sum_in(spare_reg_psum_29_11), .reg_activation(spare_reg_activation_30_11), .reg_weight(spare_reg_weight_30_11), .reg_partial_sum(spare_reg_psum_30_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_12( .activation_in(spare_reg_activation_30_11), .weight_in(spare_reg_weight_29_12), .partial_sum_in(spare_reg_psum_29_12), .reg_activation(spare_reg_activation_30_12), .reg_weight(spare_reg_weight_30_12), .reg_partial_sum(spare_reg_psum_30_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_13( .activation_in(spare_reg_activation_30_12), .weight_in(spare_reg_weight_29_13), .partial_sum_in(spare_reg_psum_29_13), .reg_activation(spare_reg_activation_30_13), .reg_weight(spare_reg_weight_30_13), .reg_partial_sum(spare_reg_psum_30_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_14( .activation_in(spare_reg_activation_30_13), .weight_in(spare_reg_weight_29_14), .partial_sum_in(spare_reg_psum_29_14), .reg_activation(spare_reg_activation_30_14), .reg_weight(spare_reg_weight_30_14), .reg_partial_sum(spare_reg_psum_30_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_15( .activation_in(spare_reg_activation_30_14), .weight_in(spare_reg_weight_29_15), .partial_sum_in(spare_reg_psum_29_15), .reg_activation(spare_reg_activation_30_15), .reg_weight(spare_reg_weight_30_15), .reg_partial_sum(spare_reg_psum_30_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_16( .activation_in(spare_reg_activation_30_15), .weight_in(spare_reg_weight_29_16), .partial_sum_in(spare_reg_psum_29_16), .reg_activation(spare_reg_activation_30_16), .reg_weight(spare_reg_weight_30_16), .reg_partial_sum(spare_reg_psum_30_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_17( .activation_in(spare_reg_activation_30_16), .weight_in(spare_reg_weight_29_17), .partial_sum_in(spare_reg_psum_29_17), .reg_activation(spare_reg_activation_30_17), .reg_weight(spare_reg_weight_30_17), .reg_partial_sum(spare_reg_psum_30_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_18( .activation_in(spare_reg_activation_30_17), .weight_in(spare_reg_weight_29_18), .partial_sum_in(spare_reg_psum_29_18), .reg_activation(spare_reg_activation_30_18), .reg_weight(spare_reg_weight_30_18), .reg_partial_sum(spare_reg_psum_30_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_19( .activation_in(spare_reg_activation_30_18), .weight_in(spare_reg_weight_29_19), .partial_sum_in(spare_reg_psum_29_19), .reg_activation(spare_reg_activation_30_19), .reg_weight(spare_reg_weight_30_19), .reg_partial_sum(spare_reg_psum_30_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_20( .activation_in(spare_reg_activation_30_19), .weight_in(spare_reg_weight_29_20), .partial_sum_in(spare_reg_psum_29_20), .reg_activation(spare_reg_activation_30_20), .reg_weight(spare_reg_weight_30_20), .reg_partial_sum(spare_reg_psum_30_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_21( .activation_in(spare_reg_activation_30_20), .weight_in(spare_reg_weight_29_21), .partial_sum_in(spare_reg_psum_29_21), .reg_activation(spare_reg_activation_30_21), .reg_weight(spare_reg_weight_30_21), .reg_partial_sum(spare_reg_psum_30_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_22( .activation_in(spare_reg_activation_30_21), .weight_in(spare_reg_weight_29_22), .partial_sum_in(spare_reg_psum_29_22), .reg_activation(spare_reg_activation_30_22), .reg_weight(spare_reg_weight_30_22), .reg_partial_sum(spare_reg_psum_30_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_23( .activation_in(spare_reg_activation_30_22), .weight_in(spare_reg_weight_29_23), .partial_sum_in(spare_reg_psum_29_23), .reg_activation(spare_reg_activation_30_23), .reg_weight(spare_reg_weight_30_23), .reg_partial_sum(spare_reg_psum_30_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_24( .activation_in(spare_reg_activation_30_23), .weight_in(spare_reg_weight_29_24), .partial_sum_in(spare_reg_psum_29_24), .reg_activation(spare_reg_activation_30_24), .reg_weight(spare_reg_weight_30_24), .reg_partial_sum(spare_reg_psum_30_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_25( .activation_in(spare_reg_activation_30_24), .weight_in(spare_reg_weight_29_25), .partial_sum_in(spare_reg_psum_29_25), .reg_activation(spare_reg_activation_30_25), .reg_weight(spare_reg_weight_30_25), .reg_partial_sum(spare_reg_psum_30_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_26( .activation_in(spare_reg_activation_30_25), .weight_in(spare_reg_weight_29_26), .partial_sum_in(spare_reg_psum_29_26), .reg_activation(spare_reg_activation_30_26), .reg_weight(spare_reg_weight_30_26), .reg_partial_sum(spare_reg_psum_30_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_27( .activation_in(spare_reg_activation_30_26), .weight_in(spare_reg_weight_29_27), .partial_sum_in(spare_reg_psum_29_27), .reg_activation(spare_reg_activation_30_27), .reg_weight(spare_reg_weight_30_27), .reg_partial_sum(spare_reg_psum_30_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_28( .activation_in(spare_reg_activation_30_27), .weight_in(spare_reg_weight_29_28), .partial_sum_in(spare_reg_psum_29_28), .reg_activation(spare_reg_activation_30_28), .reg_weight(spare_reg_weight_30_28), .reg_partial_sum(spare_reg_psum_30_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_29( .activation_in(spare_reg_activation_30_28), .weight_in(spare_reg_weight_29_29), .partial_sum_in(spare_reg_psum_29_29), .reg_activation(spare_reg_activation_30_29), .reg_weight(spare_reg_weight_30_29), .reg_partial_sum(spare_reg_psum_30_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_30( .activation_in(spare_reg_activation_30_29), .weight_in(spare_reg_weight_29_30), .partial_sum_in(spare_reg_psum_29_30), .reg_activation(spare_reg_activation_30_30), .reg_weight(spare_reg_weight_30_30), .reg_partial_sum(spare_reg_psum_30_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X30_31( .activation_in(spare_reg_activation_30_30), .weight_in(spare_reg_weight_29_31), .partial_sum_in(spare_reg_psum_29_31), .reg_weight(spare_reg_weight_30_31), .reg_partial_sum(spare_reg_psum_30_31), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_0( .activation_in(in_activation_31), .weight_in(spare_reg_weight_30_0), .partial_sum_in(spare_reg_psum_30_0), .reg_activation(spare_reg_activation_31_0), .reg_partial_sum(spare_reg_psum_31_0), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_1( .activation_in(spare_reg_activation_31_0), .weight_in(spare_reg_weight_30_1), .partial_sum_in(spare_reg_psum_30_1), .reg_activation(spare_reg_activation_31_1), .reg_partial_sum(spare_reg_psum_31_1), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_2( .activation_in(spare_reg_activation_31_1), .weight_in(spare_reg_weight_30_2), .partial_sum_in(spare_reg_psum_30_2), .reg_activation(spare_reg_activation_31_2), .reg_partial_sum(spare_reg_psum_31_2), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_3( .activation_in(spare_reg_activation_31_2), .weight_in(spare_reg_weight_30_3), .partial_sum_in(spare_reg_psum_30_3), .reg_activation(spare_reg_activation_31_3), .reg_partial_sum(spare_reg_psum_31_3), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_4( .activation_in(spare_reg_activation_31_3), .weight_in(spare_reg_weight_30_4), .partial_sum_in(spare_reg_psum_30_4), .reg_activation(spare_reg_activation_31_4), .reg_partial_sum(spare_reg_psum_31_4), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_5( .activation_in(spare_reg_activation_31_4), .weight_in(spare_reg_weight_30_5), .partial_sum_in(spare_reg_psum_30_5), .reg_activation(spare_reg_activation_31_5), .reg_partial_sum(spare_reg_psum_31_5), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_6( .activation_in(spare_reg_activation_31_5), .weight_in(spare_reg_weight_30_6), .partial_sum_in(spare_reg_psum_30_6), .reg_activation(spare_reg_activation_31_6), .reg_partial_sum(spare_reg_psum_31_6), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_7( .activation_in(spare_reg_activation_31_6), .weight_in(spare_reg_weight_30_7), .partial_sum_in(spare_reg_psum_30_7), .reg_activation(spare_reg_activation_31_7), .reg_partial_sum(spare_reg_psum_31_7), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_8( .activation_in(spare_reg_activation_31_7), .weight_in(spare_reg_weight_30_8), .partial_sum_in(spare_reg_psum_30_8), .reg_activation(spare_reg_activation_31_8), .reg_partial_sum(spare_reg_psum_31_8), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_9( .activation_in(spare_reg_activation_31_8), .weight_in(spare_reg_weight_30_9), .partial_sum_in(spare_reg_psum_30_9), .reg_activation(spare_reg_activation_31_9), .reg_partial_sum(spare_reg_psum_31_9), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_10( .activation_in(spare_reg_activation_31_9), .weight_in(spare_reg_weight_30_10), .partial_sum_in(spare_reg_psum_30_10), .reg_activation(spare_reg_activation_31_10), .reg_partial_sum(spare_reg_psum_31_10), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_11( .activation_in(spare_reg_activation_31_10), .weight_in(spare_reg_weight_30_11), .partial_sum_in(spare_reg_psum_30_11), .reg_activation(spare_reg_activation_31_11), .reg_partial_sum(spare_reg_psum_31_11), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_12( .activation_in(spare_reg_activation_31_11), .weight_in(spare_reg_weight_30_12), .partial_sum_in(spare_reg_psum_30_12), .reg_activation(spare_reg_activation_31_12), .reg_partial_sum(spare_reg_psum_31_12), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_13( .activation_in(spare_reg_activation_31_12), .weight_in(spare_reg_weight_30_13), .partial_sum_in(spare_reg_psum_30_13), .reg_activation(spare_reg_activation_31_13), .reg_partial_sum(spare_reg_psum_31_13), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_14( .activation_in(spare_reg_activation_31_13), .weight_in(spare_reg_weight_30_14), .partial_sum_in(spare_reg_psum_30_14), .reg_activation(spare_reg_activation_31_14), .reg_partial_sum(spare_reg_psum_31_14), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_15( .activation_in(spare_reg_activation_31_14), .weight_in(spare_reg_weight_30_15), .partial_sum_in(spare_reg_psum_30_15), .reg_activation(spare_reg_activation_31_15), .reg_partial_sum(spare_reg_psum_31_15), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_16( .activation_in(spare_reg_activation_31_15), .weight_in(spare_reg_weight_30_16), .partial_sum_in(spare_reg_psum_30_16), .reg_activation(spare_reg_activation_31_16), .reg_partial_sum(spare_reg_psum_31_16), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_17( .activation_in(spare_reg_activation_31_16), .weight_in(spare_reg_weight_30_17), .partial_sum_in(spare_reg_psum_30_17), .reg_activation(spare_reg_activation_31_17), .reg_partial_sum(spare_reg_psum_31_17), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_18( .activation_in(spare_reg_activation_31_17), .weight_in(spare_reg_weight_30_18), .partial_sum_in(spare_reg_psum_30_18), .reg_activation(spare_reg_activation_31_18), .reg_partial_sum(spare_reg_psum_31_18), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_19( .activation_in(spare_reg_activation_31_18), .weight_in(spare_reg_weight_30_19), .partial_sum_in(spare_reg_psum_30_19), .reg_activation(spare_reg_activation_31_19), .reg_partial_sum(spare_reg_psum_31_19), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_20( .activation_in(spare_reg_activation_31_19), .weight_in(spare_reg_weight_30_20), .partial_sum_in(spare_reg_psum_30_20), .reg_activation(spare_reg_activation_31_20), .reg_partial_sum(spare_reg_psum_31_20), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_21( .activation_in(spare_reg_activation_31_20), .weight_in(spare_reg_weight_30_21), .partial_sum_in(spare_reg_psum_30_21), .reg_activation(spare_reg_activation_31_21), .reg_partial_sum(spare_reg_psum_31_21), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_22( .activation_in(spare_reg_activation_31_21), .weight_in(spare_reg_weight_30_22), .partial_sum_in(spare_reg_psum_30_22), .reg_activation(spare_reg_activation_31_22), .reg_partial_sum(spare_reg_psum_31_22), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_23( .activation_in(spare_reg_activation_31_22), .weight_in(spare_reg_weight_30_23), .partial_sum_in(spare_reg_psum_30_23), .reg_activation(spare_reg_activation_31_23), .reg_partial_sum(spare_reg_psum_31_23), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_24( .activation_in(spare_reg_activation_31_23), .weight_in(spare_reg_weight_30_24), .partial_sum_in(spare_reg_psum_30_24), .reg_activation(spare_reg_activation_31_24), .reg_partial_sum(spare_reg_psum_31_24), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_25( .activation_in(spare_reg_activation_31_24), .weight_in(spare_reg_weight_30_25), .partial_sum_in(spare_reg_psum_30_25), .reg_activation(spare_reg_activation_31_25), .reg_partial_sum(spare_reg_psum_31_25), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_26( .activation_in(spare_reg_activation_31_25), .weight_in(spare_reg_weight_30_26), .partial_sum_in(spare_reg_psum_30_26), .reg_activation(spare_reg_activation_31_26), .reg_partial_sum(spare_reg_psum_31_26), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_27( .activation_in(spare_reg_activation_31_26), .weight_in(spare_reg_weight_30_27), .partial_sum_in(spare_reg_psum_30_27), .reg_activation(spare_reg_activation_31_27), .reg_partial_sum(spare_reg_psum_31_27), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_28( .activation_in(spare_reg_activation_31_27), .weight_in(spare_reg_weight_30_28), .partial_sum_in(spare_reg_psum_30_28), .reg_activation(spare_reg_activation_31_28), .reg_partial_sum(spare_reg_psum_31_28), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_29( .activation_in(spare_reg_activation_31_28), .weight_in(spare_reg_weight_30_29), .partial_sum_in(spare_reg_psum_30_29), .reg_activation(spare_reg_activation_31_29), .reg_partial_sum(spare_reg_psum_31_29), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_30( .activation_in(spare_reg_activation_31_29), .weight_in(spare_reg_weight_30_30), .partial_sum_in(spare_reg_psum_30_30), .reg_activation(spare_reg_activation_31_30), .reg_partial_sum(spare_reg_psum_31_30), .clk(clk), .rst(rst), .weight_en(weight_en));
PE X31_31( .activation_in(spare_reg_activation_31_30), .weight_in(spare_reg_weight_30_31), .partial_sum_in(spare_reg_psum_30_31), .reg_partial_sum(spare_reg_psum_31_31), .clk(clk), .rst(rst), .weight_en(weight_en));
endmodule