`include "/home/wzc/verilog/systolic_array/SA22.v"
module SA64(rst, clk, weight_en, in_weight1_1_1, in_psum1_1_1, in_weight1_1_2, in_psum1_1_2, in_weight1_2_1, in_psum1_2_1, in_weight1_2_2, in_psum1_2_2, in_weight1_3_1, in_psum1_3_1, in_weight1_3_2, in_psum1_3_2, in_weight1_4_1, in_psum1_4_1, in_weight1_4_2, in_psum1_4_2, in_weight1_5_1, in_psum1_5_1, in_weight1_5_2, in_psum1_5_2, in_weight1_6_1, in_psum1_6_1, in_weight1_6_2, in_psum1_6_2, in_weight1_7_1, in_psum1_7_1, in_weight1_7_2, in_psum1_7_2, in_weight1_8_1, in_psum1_8_1, in_weight1_8_2, in_psum1_8_2, in_weight1_9_1, in_psum1_9_1, in_weight1_9_2, in_psum1_9_2, in_weight1_10_1, in_psum1_10_1, in_weight1_10_2, in_psum1_10_2, in_weight1_11_1, in_psum1_11_1, in_weight1_11_2, in_psum1_11_2, in_weight1_12_1, in_psum1_12_1, in_weight1_12_2, in_psum1_12_2, in_weight1_13_1, in_psum1_13_1, in_weight1_13_2, in_psum1_13_2, in_weight1_14_1, in_psum1_14_1, in_weight1_14_2, in_psum1_14_2, in_weight1_15_1, in_psum1_15_1, in_weight1_15_2, in_psum1_15_2, in_weight1_16_1, in_psum1_16_1, in_weight1_16_2, in_psum1_16_2, in_weight1_17_1, in_psum1_17_1, in_weight1_17_2, in_psum1_17_2, in_weight1_18_1, in_psum1_18_1, in_weight1_18_2, in_psum1_18_2, in_weight1_19_1, in_psum1_19_1, in_weight1_19_2, in_psum1_19_2, in_weight1_20_1, in_psum1_20_1, in_weight1_20_2, in_psum1_20_2, in_weight1_21_1, in_psum1_21_1, in_weight1_21_2, in_psum1_21_2, in_weight1_22_1, in_psum1_22_1, in_weight1_22_2, in_psum1_22_2, in_weight1_23_1, in_psum1_23_1, in_weight1_23_2, in_psum1_23_2, in_weight1_24_1, in_psum1_24_1, in_weight1_24_2, in_psum1_24_2, in_weight1_25_1, in_psum1_25_1, in_weight1_25_2, in_psum1_25_2, in_weight1_26_1, in_psum1_26_1, in_weight1_26_2, in_psum1_26_2, in_weight1_27_1, in_psum1_27_1, in_weight1_27_2, in_psum1_27_2, in_weight1_28_1, in_psum1_28_1, in_weight1_28_2, in_psum1_28_2, in_weight1_29_1, in_psum1_29_1, in_weight1_29_2, in_psum1_29_2, in_weight1_30_1, in_psum1_30_1, in_weight1_30_2, in_psum1_30_2, in_weight1_31_1, in_psum1_31_1, in_weight1_31_2, in_psum1_31_2, in_weight1_32_1, in_psum1_32_1, in_weight1_32_2, in_psum1_32_2, in_activation1_1_1, in_activation1_1_2, in_activation2_1_1, in_activation2_1_2, in_activation3_1_1, in_activation3_1_2, in_activation4_1_1, in_activation4_1_2, in_activation5_1_1, in_activation5_1_2, in_activation6_1_1, in_activation6_1_2, in_activation7_1_1, in_activation7_1_2, in_activation8_1_1, in_activation8_1_2, in_activation9_1_1, in_activation9_1_2, in_activation10_1_1, in_activation10_1_2, in_activation11_1_1, in_activation11_1_2, in_activation12_1_1, in_activation12_1_2, in_activation13_1_1, in_activation13_1_2, in_activation14_1_1, in_activation14_1_2, in_activation15_1_1, in_activation15_1_2, in_activation16_1_1, in_activation16_1_2, in_activation17_1_1, in_activation17_1_2, in_activation18_1_1, in_activation18_1_2, in_activation19_1_1, in_activation19_1_2, in_activation20_1_1, in_activation20_1_2, in_activation21_1_1, in_activation21_1_2, in_activation22_1_1, in_activation22_1_2, in_activation23_1_1, in_activation23_1_2, in_activation24_1_1, in_activation24_1_2, in_activation25_1_1, in_activation25_1_2, in_activation26_1_1, in_activation26_1_2, in_activation27_1_1, in_activation27_1_2, in_activation28_1_1, in_activation28_1_2, in_activation29_1_1, in_activation29_1_2, in_activation30_1_1, in_activation30_1_2, in_activation31_1_1, in_activation31_1_2, in_activation32_1_1, in_activation32_1_2, reg_psum32_1_1, reg_psum32_1_2, reg_psum32_2_1, reg_psum32_2_2, reg_psum32_3_1, reg_psum32_3_2, reg_psum32_4_1, reg_psum32_4_2, reg_psum32_5_1, reg_psum32_5_2, reg_psum32_6_1, reg_psum32_6_2, reg_psum32_7_1, reg_psum32_7_2, reg_psum32_8_1, reg_psum32_8_2, reg_psum32_9_1, reg_psum32_9_2, reg_psum32_10_1, reg_psum32_10_2, reg_psum32_11_1, reg_psum32_11_2, reg_psum32_12_1, reg_psum32_12_2, reg_psum32_13_1, reg_psum32_13_2, reg_psum32_14_1, reg_psum32_14_2, reg_psum32_15_1, reg_psum32_15_2, reg_psum32_16_1, reg_psum32_16_2, reg_psum32_17_1, reg_psum32_17_2, reg_psum32_18_1, reg_psum32_18_2, reg_psum32_19_1, reg_psum32_19_2, reg_psum32_20_1, reg_psum32_20_2, reg_psum32_21_1, reg_psum32_21_2, reg_psum32_22_1, reg_psum32_22_2, reg_psum32_23_1, reg_psum32_23_2, reg_psum32_24_1, reg_psum32_24_2, reg_psum32_25_1, reg_psum32_25_2, reg_psum32_26_1, reg_psum32_26_2, reg_psum32_27_1, reg_psum32_27_2, reg_psum32_28_1, reg_psum32_28_2, reg_psum32_29_1, reg_psum32_29_2, reg_psum32_30_1, reg_psum32_30_2, reg_psum32_31_1, reg_psum32_31_2, reg_psum32_32_1, reg_psum32_32_2);

input weight_en;
input clk,rst;
input[15:0]   in_weight1_1_1;
input[15:0]   in_psum1_1_1;
input[15:0]   in_weight1_1_2;
input[15:0]   in_psum1_1_2;
input[15:0]   in_weight1_2_1;
input[15:0]   in_psum1_2_1;
input[15:0]   in_weight1_2_2;
input[15:0]   in_psum1_2_2;
input[15:0]   in_weight1_3_1;
input[15:0]   in_psum1_3_1;
input[15:0]   in_weight1_3_2;
input[15:0]   in_psum1_3_2;
input[15:0]   in_weight1_4_1;
input[15:0]   in_psum1_4_1;
input[15:0]   in_weight1_4_2;
input[15:0]   in_psum1_4_2;
input[15:0]   in_weight1_5_1;
input[15:0]   in_psum1_5_1;
input[15:0]   in_weight1_5_2;
input[15:0]   in_psum1_5_2;
input[15:0]   in_weight1_6_1;
input[15:0]   in_psum1_6_1;
input[15:0]   in_weight1_6_2;
input[15:0]   in_psum1_6_2;
input[15:0]   in_weight1_7_1;
input[15:0]   in_psum1_7_1;
input[15:0]   in_weight1_7_2;
input[15:0]   in_psum1_7_2;
input[15:0]   in_weight1_8_1;
input[15:0]   in_psum1_8_1;
input[15:0]   in_weight1_8_2;
input[15:0]   in_psum1_8_2;
input[15:0]   in_weight1_9_1;
input[15:0]   in_psum1_9_1;
input[15:0]   in_weight1_9_2;
input[15:0]   in_psum1_9_2;
input[15:0]   in_weight1_10_1;
input[15:0]   in_psum1_10_1;
input[15:0]   in_weight1_10_2;
input[15:0]   in_psum1_10_2;
input[15:0]   in_weight1_11_1;
input[15:0]   in_psum1_11_1;
input[15:0]   in_weight1_11_2;
input[15:0]   in_psum1_11_2;
input[15:0]   in_weight1_12_1;
input[15:0]   in_psum1_12_1;
input[15:0]   in_weight1_12_2;
input[15:0]   in_psum1_12_2;
input[15:0]   in_weight1_13_1;
input[15:0]   in_psum1_13_1;
input[15:0]   in_weight1_13_2;
input[15:0]   in_psum1_13_2;
input[15:0]   in_weight1_14_1;
input[15:0]   in_psum1_14_1;
input[15:0]   in_weight1_14_2;
input[15:0]   in_psum1_14_2;
input[15:0]   in_weight1_15_1;
input[15:0]   in_psum1_15_1;
input[15:0]   in_weight1_15_2;
input[15:0]   in_psum1_15_2;
input[15:0]   in_weight1_16_1;
input[15:0]   in_psum1_16_1;
input[15:0]   in_weight1_16_2;
input[15:0]   in_psum1_16_2;
input[15:0]   in_weight1_17_1;
input[15:0]   in_psum1_17_1;
input[15:0]   in_weight1_17_2;
input[15:0]   in_psum1_17_2;
input[15:0]   in_weight1_18_1;
input[15:0]   in_psum1_18_1;
input[15:0]   in_weight1_18_2;
input[15:0]   in_psum1_18_2;
input[15:0]   in_weight1_19_1;
input[15:0]   in_psum1_19_1;
input[15:0]   in_weight1_19_2;
input[15:0]   in_psum1_19_2;
input[15:0]   in_weight1_20_1;
input[15:0]   in_psum1_20_1;
input[15:0]   in_weight1_20_2;
input[15:0]   in_psum1_20_2;
input[15:0]   in_weight1_21_1;
input[15:0]   in_psum1_21_1;
input[15:0]   in_weight1_21_2;
input[15:0]   in_psum1_21_2;
input[15:0]   in_weight1_22_1;
input[15:0]   in_psum1_22_1;
input[15:0]   in_weight1_22_2;
input[15:0]   in_psum1_22_2;
input[15:0]   in_weight1_23_1;
input[15:0]   in_psum1_23_1;
input[15:0]   in_weight1_23_2;
input[15:0]   in_psum1_23_2;
input[15:0]   in_weight1_24_1;
input[15:0]   in_psum1_24_1;
input[15:0]   in_weight1_24_2;
input[15:0]   in_psum1_24_2;
input[15:0]   in_weight1_25_1;
input[15:0]   in_psum1_25_1;
input[15:0]   in_weight1_25_2;
input[15:0]   in_psum1_25_2;
input[15:0]   in_weight1_26_1;
input[15:0]   in_psum1_26_1;
input[15:0]   in_weight1_26_2;
input[15:0]   in_psum1_26_2;
input[15:0]   in_weight1_27_1;
input[15:0]   in_psum1_27_1;
input[15:0]   in_weight1_27_2;
input[15:0]   in_psum1_27_2;
input[15:0]   in_weight1_28_1;
input[15:0]   in_psum1_28_1;
input[15:0]   in_weight1_28_2;
input[15:0]   in_psum1_28_2;
input[15:0]   in_weight1_29_1;
input[15:0]   in_psum1_29_1;
input[15:0]   in_weight1_29_2;
input[15:0]   in_psum1_29_2;
input[15:0]   in_weight1_30_1;
input[15:0]   in_psum1_30_1;
input[15:0]   in_weight1_30_2;
input[15:0]   in_psum1_30_2;
input[15:0]   in_weight1_31_1;
input[15:0]   in_psum1_31_1;
input[15:0]   in_weight1_31_2;
input[15:0]   in_psum1_31_2;
input[15:0]   in_weight1_32_1;
input[15:0]   in_psum1_32_1;
input[15:0]   in_weight1_32_2;
input[15:0]   in_psum1_32_2;
input[15:0]   in_activation1_1_1;
input[15:0]   in_activation1_1_2;
input[15:0]   in_activation2_1_1;
input[15:0]   in_activation2_1_2;
input[15:0]   in_activation3_1_1;
input[15:0]   in_activation3_1_2;
input[15:0]   in_activation4_1_1;
input[15:0]   in_activation4_1_2;
input[15:0]   in_activation5_1_1;
input[15:0]   in_activation5_1_2;
input[15:0]   in_activation6_1_1;
input[15:0]   in_activation6_1_2;
input[15:0]   in_activation7_1_1;
input[15:0]   in_activation7_1_2;
input[15:0]   in_activation8_1_1;
input[15:0]   in_activation8_1_2;
input[15:0]   in_activation9_1_1;
input[15:0]   in_activation9_1_2;
input[15:0]   in_activation10_1_1;
input[15:0]   in_activation10_1_2;
input[15:0]   in_activation11_1_1;
input[15:0]   in_activation11_1_2;
input[15:0]   in_activation12_1_1;
input[15:0]   in_activation12_1_2;
input[15:0]   in_activation13_1_1;
input[15:0]   in_activation13_1_2;
input[15:0]   in_activation14_1_1;
input[15:0]   in_activation14_1_2;
input[15:0]   in_activation15_1_1;
input[15:0]   in_activation15_1_2;
input[15:0]   in_activation16_1_1;
input[15:0]   in_activation16_1_2;
input[15:0]   in_activation17_1_1;
input[15:0]   in_activation17_1_2;
input[15:0]   in_activation18_1_1;
input[15:0]   in_activation18_1_2;
input[15:0]   in_activation19_1_1;
input[15:0]   in_activation19_1_2;
input[15:0]   in_activation20_1_1;
input[15:0]   in_activation20_1_2;
input[15:0]   in_activation21_1_1;
input[15:0]   in_activation21_1_2;
input[15:0]   in_activation22_1_1;
input[15:0]   in_activation22_1_2;
input[15:0]   in_activation23_1_1;
input[15:0]   in_activation23_1_2;
input[15:0]   in_activation24_1_1;
input[15:0]   in_activation24_1_2;
input[15:0]   in_activation25_1_1;
input[15:0]   in_activation25_1_2;
input[15:0]   in_activation26_1_1;
input[15:0]   in_activation26_1_2;
input[15:0]   in_activation27_1_1;
input[15:0]   in_activation27_1_2;
input[15:0]   in_activation28_1_1;
input[15:0]   in_activation28_1_2;
input[15:0]   in_activation29_1_1;
input[15:0]   in_activation29_1_2;
input[15:0]   in_activation30_1_1;
input[15:0]   in_activation30_1_2;
input[15:0]   in_activation31_1_1;
input[15:0]   in_activation31_1_2;
input[15:0]   in_activation32_1_1;
input[15:0]   in_activation32_1_2;
output[15:0]   reg_psum32_1_1;
output[15:0]   reg_psum32_1_2;
output[15:0]   reg_psum32_2_1;
output[15:0]   reg_psum32_2_2;
output[15:0]   reg_psum32_3_1;
output[15:0]   reg_psum32_3_2;
output[15:0]   reg_psum32_4_1;
output[15:0]   reg_psum32_4_2;
output[15:0]   reg_psum32_5_1;
output[15:0]   reg_psum32_5_2;
output[15:0]   reg_psum32_6_1;
output[15:0]   reg_psum32_6_2;
output[15:0]   reg_psum32_7_1;
output[15:0]   reg_psum32_7_2;
output[15:0]   reg_psum32_8_1;
output[15:0]   reg_psum32_8_2;
output[15:0]   reg_psum32_9_1;
output[15:0]   reg_psum32_9_2;
output[15:0]   reg_psum32_10_1;
output[15:0]   reg_psum32_10_2;
output[15:0]   reg_psum32_11_1;
output[15:0]   reg_psum32_11_2;
output[15:0]   reg_psum32_12_1;
output[15:0]   reg_psum32_12_2;
output[15:0]   reg_psum32_13_1;
output[15:0]   reg_psum32_13_2;
output[15:0]   reg_psum32_14_1;
output[15:0]   reg_psum32_14_2;
output[15:0]   reg_psum32_15_1;
output[15:0]   reg_psum32_15_2;
output[15:0]   reg_psum32_16_1;
output[15:0]   reg_psum32_16_2;
output[15:0]   reg_psum32_17_1;
output[15:0]   reg_psum32_17_2;
output[15:0]   reg_psum32_18_1;
output[15:0]   reg_psum32_18_2;
output[15:0]   reg_psum32_19_1;
output[15:0]   reg_psum32_19_2;
output[15:0]   reg_psum32_20_1;
output[15:0]   reg_psum32_20_2;
output[15:0]   reg_psum32_21_1;
output[15:0]   reg_psum32_21_2;
output[15:0]   reg_psum32_22_1;
output[15:0]   reg_psum32_22_2;
output[15:0]   reg_psum32_23_1;
output[15:0]   reg_psum32_23_2;
output[15:0]   reg_psum32_24_1;
output[15:0]   reg_psum32_24_2;
output[15:0]   reg_psum32_25_1;
output[15:0]   reg_psum32_25_2;
output[15:0]   reg_psum32_26_1;
output[15:0]   reg_psum32_26_2;
output[15:0]   reg_psum32_27_1;
output[15:0]   reg_psum32_27_2;
output[15:0]   reg_psum32_28_1;
output[15:0]   reg_psum32_28_2;
output[15:0]   reg_psum32_29_1;
output[15:0]   reg_psum32_29_2;
output[15:0]   reg_psum32_30_1;
output[15:0]   reg_psum32_30_2;
output[15:0]   reg_psum32_31_1;
output[15:0]   reg_psum32_31_2;
output[15:0]   reg_psum32_32_1;
output[15:0]   reg_psum32_32_2;
wire[15:0]    reg_activation1_1_1;
wire[15:0]    reg_activation1_1_2;
wire[15:0]    reg_activation1_2_1;
wire[15:0]    reg_activation1_2_2;
wire[15:0]    reg_activation1_3_1;
wire[15:0]    reg_activation1_3_2;
wire[15:0]    reg_activation1_4_1;
wire[15:0]    reg_activation1_4_2;
wire[15:0]    reg_activation1_5_1;
wire[15:0]    reg_activation1_5_2;
wire[15:0]    reg_activation1_6_1;
wire[15:0]    reg_activation1_6_2;
wire[15:0]    reg_activation1_7_1;
wire[15:0]    reg_activation1_7_2;
wire[15:0]    reg_activation1_8_1;
wire[15:0]    reg_activation1_8_2;
wire[15:0]    reg_activation1_9_1;
wire[15:0]    reg_activation1_9_2;
wire[15:0]    reg_activation1_10_1;
wire[15:0]    reg_activation1_10_2;
wire[15:0]    reg_activation1_11_1;
wire[15:0]    reg_activation1_11_2;
wire[15:0]    reg_activation1_12_1;
wire[15:0]    reg_activation1_12_2;
wire[15:0]    reg_activation1_13_1;
wire[15:0]    reg_activation1_13_2;
wire[15:0]    reg_activation1_14_1;
wire[15:0]    reg_activation1_14_2;
wire[15:0]    reg_activation1_15_1;
wire[15:0]    reg_activation1_15_2;
wire[15:0]    reg_activation1_16_1;
wire[15:0]    reg_activation1_16_2;
wire[15:0]    reg_activation1_17_1;
wire[15:0]    reg_activation1_17_2;
wire[15:0]    reg_activation1_18_1;
wire[15:0]    reg_activation1_18_2;
wire[15:0]    reg_activation1_19_1;
wire[15:0]    reg_activation1_19_2;
wire[15:0]    reg_activation1_20_1;
wire[15:0]    reg_activation1_20_2;
wire[15:0]    reg_activation1_21_1;
wire[15:0]    reg_activation1_21_2;
wire[15:0]    reg_activation1_22_1;
wire[15:0]    reg_activation1_22_2;
wire[15:0]    reg_activation1_23_1;
wire[15:0]    reg_activation1_23_2;
wire[15:0]    reg_activation1_24_1;
wire[15:0]    reg_activation1_24_2;
wire[15:0]    reg_activation1_25_1;
wire[15:0]    reg_activation1_25_2;
wire[15:0]    reg_activation1_26_1;
wire[15:0]    reg_activation1_26_2;
wire[15:0]    reg_activation1_27_1;
wire[15:0]    reg_activation1_27_2;
wire[15:0]    reg_activation1_28_1;
wire[15:0]    reg_activation1_28_2;
wire[15:0]    reg_activation1_29_1;
wire[15:0]    reg_activation1_29_2;
wire[15:0]    reg_activation1_30_1;
wire[15:0]    reg_activation1_30_2;
wire[15:0]    reg_activation1_31_1;
wire[15:0]    reg_activation1_31_2;
wire[15:0]    reg_activation2_1_1;
wire[15:0]    reg_activation2_1_2;
wire[15:0]    reg_activation2_2_1;
wire[15:0]    reg_activation2_2_2;
wire[15:0]    reg_activation2_3_1;
wire[15:0]    reg_activation2_3_2;
wire[15:0]    reg_activation2_4_1;
wire[15:0]    reg_activation2_4_2;
wire[15:0]    reg_activation2_5_1;
wire[15:0]    reg_activation2_5_2;
wire[15:0]    reg_activation2_6_1;
wire[15:0]    reg_activation2_6_2;
wire[15:0]    reg_activation2_7_1;
wire[15:0]    reg_activation2_7_2;
wire[15:0]    reg_activation2_8_1;
wire[15:0]    reg_activation2_8_2;
wire[15:0]    reg_activation2_9_1;
wire[15:0]    reg_activation2_9_2;
wire[15:0]    reg_activation2_10_1;
wire[15:0]    reg_activation2_10_2;
wire[15:0]    reg_activation2_11_1;
wire[15:0]    reg_activation2_11_2;
wire[15:0]    reg_activation2_12_1;
wire[15:0]    reg_activation2_12_2;
wire[15:0]    reg_activation2_13_1;
wire[15:0]    reg_activation2_13_2;
wire[15:0]    reg_activation2_14_1;
wire[15:0]    reg_activation2_14_2;
wire[15:0]    reg_activation2_15_1;
wire[15:0]    reg_activation2_15_2;
wire[15:0]    reg_activation2_16_1;
wire[15:0]    reg_activation2_16_2;
wire[15:0]    reg_activation2_17_1;
wire[15:0]    reg_activation2_17_2;
wire[15:0]    reg_activation2_18_1;
wire[15:0]    reg_activation2_18_2;
wire[15:0]    reg_activation2_19_1;
wire[15:0]    reg_activation2_19_2;
wire[15:0]    reg_activation2_20_1;
wire[15:0]    reg_activation2_20_2;
wire[15:0]    reg_activation2_21_1;
wire[15:0]    reg_activation2_21_2;
wire[15:0]    reg_activation2_22_1;
wire[15:0]    reg_activation2_22_2;
wire[15:0]    reg_activation2_23_1;
wire[15:0]    reg_activation2_23_2;
wire[15:0]    reg_activation2_24_1;
wire[15:0]    reg_activation2_24_2;
wire[15:0]    reg_activation2_25_1;
wire[15:0]    reg_activation2_25_2;
wire[15:0]    reg_activation2_26_1;
wire[15:0]    reg_activation2_26_2;
wire[15:0]    reg_activation2_27_1;
wire[15:0]    reg_activation2_27_2;
wire[15:0]    reg_activation2_28_1;
wire[15:0]    reg_activation2_28_2;
wire[15:0]    reg_activation2_29_1;
wire[15:0]    reg_activation2_29_2;
wire[15:0]    reg_activation2_30_1;
wire[15:0]    reg_activation2_30_2;
wire[15:0]    reg_activation2_31_1;
wire[15:0]    reg_activation2_31_2;
wire[15:0]    reg_activation3_1_1;
wire[15:0]    reg_activation3_1_2;
wire[15:0]    reg_activation3_2_1;
wire[15:0]    reg_activation3_2_2;
wire[15:0]    reg_activation3_3_1;
wire[15:0]    reg_activation3_3_2;
wire[15:0]    reg_activation3_4_1;
wire[15:0]    reg_activation3_4_2;
wire[15:0]    reg_activation3_5_1;
wire[15:0]    reg_activation3_5_2;
wire[15:0]    reg_activation3_6_1;
wire[15:0]    reg_activation3_6_2;
wire[15:0]    reg_activation3_7_1;
wire[15:0]    reg_activation3_7_2;
wire[15:0]    reg_activation3_8_1;
wire[15:0]    reg_activation3_8_2;
wire[15:0]    reg_activation3_9_1;
wire[15:0]    reg_activation3_9_2;
wire[15:0]    reg_activation3_10_1;
wire[15:0]    reg_activation3_10_2;
wire[15:0]    reg_activation3_11_1;
wire[15:0]    reg_activation3_11_2;
wire[15:0]    reg_activation3_12_1;
wire[15:0]    reg_activation3_12_2;
wire[15:0]    reg_activation3_13_1;
wire[15:0]    reg_activation3_13_2;
wire[15:0]    reg_activation3_14_1;
wire[15:0]    reg_activation3_14_2;
wire[15:0]    reg_activation3_15_1;
wire[15:0]    reg_activation3_15_2;
wire[15:0]    reg_activation3_16_1;
wire[15:0]    reg_activation3_16_2;
wire[15:0]    reg_activation3_17_1;
wire[15:0]    reg_activation3_17_2;
wire[15:0]    reg_activation3_18_1;
wire[15:0]    reg_activation3_18_2;
wire[15:0]    reg_activation3_19_1;
wire[15:0]    reg_activation3_19_2;
wire[15:0]    reg_activation3_20_1;
wire[15:0]    reg_activation3_20_2;
wire[15:0]    reg_activation3_21_1;
wire[15:0]    reg_activation3_21_2;
wire[15:0]    reg_activation3_22_1;
wire[15:0]    reg_activation3_22_2;
wire[15:0]    reg_activation3_23_1;
wire[15:0]    reg_activation3_23_2;
wire[15:0]    reg_activation3_24_1;
wire[15:0]    reg_activation3_24_2;
wire[15:0]    reg_activation3_25_1;
wire[15:0]    reg_activation3_25_2;
wire[15:0]    reg_activation3_26_1;
wire[15:0]    reg_activation3_26_2;
wire[15:0]    reg_activation3_27_1;
wire[15:0]    reg_activation3_27_2;
wire[15:0]    reg_activation3_28_1;
wire[15:0]    reg_activation3_28_2;
wire[15:0]    reg_activation3_29_1;
wire[15:0]    reg_activation3_29_2;
wire[15:0]    reg_activation3_30_1;
wire[15:0]    reg_activation3_30_2;
wire[15:0]    reg_activation3_31_1;
wire[15:0]    reg_activation3_31_2;
wire[15:0]    reg_activation4_1_1;
wire[15:0]    reg_activation4_1_2;
wire[15:0]    reg_activation4_2_1;
wire[15:0]    reg_activation4_2_2;
wire[15:0]    reg_activation4_3_1;
wire[15:0]    reg_activation4_3_2;
wire[15:0]    reg_activation4_4_1;
wire[15:0]    reg_activation4_4_2;
wire[15:0]    reg_activation4_5_1;
wire[15:0]    reg_activation4_5_2;
wire[15:0]    reg_activation4_6_1;
wire[15:0]    reg_activation4_6_2;
wire[15:0]    reg_activation4_7_1;
wire[15:0]    reg_activation4_7_2;
wire[15:0]    reg_activation4_8_1;
wire[15:0]    reg_activation4_8_2;
wire[15:0]    reg_activation4_9_1;
wire[15:0]    reg_activation4_9_2;
wire[15:0]    reg_activation4_10_1;
wire[15:0]    reg_activation4_10_2;
wire[15:0]    reg_activation4_11_1;
wire[15:0]    reg_activation4_11_2;
wire[15:0]    reg_activation4_12_1;
wire[15:0]    reg_activation4_12_2;
wire[15:0]    reg_activation4_13_1;
wire[15:0]    reg_activation4_13_2;
wire[15:0]    reg_activation4_14_1;
wire[15:0]    reg_activation4_14_2;
wire[15:0]    reg_activation4_15_1;
wire[15:0]    reg_activation4_15_2;
wire[15:0]    reg_activation4_16_1;
wire[15:0]    reg_activation4_16_2;
wire[15:0]    reg_activation4_17_1;
wire[15:0]    reg_activation4_17_2;
wire[15:0]    reg_activation4_18_1;
wire[15:0]    reg_activation4_18_2;
wire[15:0]    reg_activation4_19_1;
wire[15:0]    reg_activation4_19_2;
wire[15:0]    reg_activation4_20_1;
wire[15:0]    reg_activation4_20_2;
wire[15:0]    reg_activation4_21_1;
wire[15:0]    reg_activation4_21_2;
wire[15:0]    reg_activation4_22_1;
wire[15:0]    reg_activation4_22_2;
wire[15:0]    reg_activation4_23_1;
wire[15:0]    reg_activation4_23_2;
wire[15:0]    reg_activation4_24_1;
wire[15:0]    reg_activation4_24_2;
wire[15:0]    reg_activation4_25_1;
wire[15:0]    reg_activation4_25_2;
wire[15:0]    reg_activation4_26_1;
wire[15:0]    reg_activation4_26_2;
wire[15:0]    reg_activation4_27_1;
wire[15:0]    reg_activation4_27_2;
wire[15:0]    reg_activation4_28_1;
wire[15:0]    reg_activation4_28_2;
wire[15:0]    reg_activation4_29_1;
wire[15:0]    reg_activation4_29_2;
wire[15:0]    reg_activation4_30_1;
wire[15:0]    reg_activation4_30_2;
wire[15:0]    reg_activation4_31_1;
wire[15:0]    reg_activation4_31_2;
wire[15:0]    reg_activation5_1_1;
wire[15:0]    reg_activation5_1_2;
wire[15:0]    reg_activation5_2_1;
wire[15:0]    reg_activation5_2_2;
wire[15:0]    reg_activation5_3_1;
wire[15:0]    reg_activation5_3_2;
wire[15:0]    reg_activation5_4_1;
wire[15:0]    reg_activation5_4_2;
wire[15:0]    reg_activation5_5_1;
wire[15:0]    reg_activation5_5_2;
wire[15:0]    reg_activation5_6_1;
wire[15:0]    reg_activation5_6_2;
wire[15:0]    reg_activation5_7_1;
wire[15:0]    reg_activation5_7_2;
wire[15:0]    reg_activation5_8_1;
wire[15:0]    reg_activation5_8_2;
wire[15:0]    reg_activation5_9_1;
wire[15:0]    reg_activation5_9_2;
wire[15:0]    reg_activation5_10_1;
wire[15:0]    reg_activation5_10_2;
wire[15:0]    reg_activation5_11_1;
wire[15:0]    reg_activation5_11_2;
wire[15:0]    reg_activation5_12_1;
wire[15:0]    reg_activation5_12_2;
wire[15:0]    reg_activation5_13_1;
wire[15:0]    reg_activation5_13_2;
wire[15:0]    reg_activation5_14_1;
wire[15:0]    reg_activation5_14_2;
wire[15:0]    reg_activation5_15_1;
wire[15:0]    reg_activation5_15_2;
wire[15:0]    reg_activation5_16_1;
wire[15:0]    reg_activation5_16_2;
wire[15:0]    reg_activation5_17_1;
wire[15:0]    reg_activation5_17_2;
wire[15:0]    reg_activation5_18_1;
wire[15:0]    reg_activation5_18_2;
wire[15:0]    reg_activation5_19_1;
wire[15:0]    reg_activation5_19_2;
wire[15:0]    reg_activation5_20_1;
wire[15:0]    reg_activation5_20_2;
wire[15:0]    reg_activation5_21_1;
wire[15:0]    reg_activation5_21_2;
wire[15:0]    reg_activation5_22_1;
wire[15:0]    reg_activation5_22_2;
wire[15:0]    reg_activation5_23_1;
wire[15:0]    reg_activation5_23_2;
wire[15:0]    reg_activation5_24_1;
wire[15:0]    reg_activation5_24_2;
wire[15:0]    reg_activation5_25_1;
wire[15:0]    reg_activation5_25_2;
wire[15:0]    reg_activation5_26_1;
wire[15:0]    reg_activation5_26_2;
wire[15:0]    reg_activation5_27_1;
wire[15:0]    reg_activation5_27_2;
wire[15:0]    reg_activation5_28_1;
wire[15:0]    reg_activation5_28_2;
wire[15:0]    reg_activation5_29_1;
wire[15:0]    reg_activation5_29_2;
wire[15:0]    reg_activation5_30_1;
wire[15:0]    reg_activation5_30_2;
wire[15:0]    reg_activation5_31_1;
wire[15:0]    reg_activation5_31_2;
wire[15:0]    reg_activation6_1_1;
wire[15:0]    reg_activation6_1_2;
wire[15:0]    reg_activation6_2_1;
wire[15:0]    reg_activation6_2_2;
wire[15:0]    reg_activation6_3_1;
wire[15:0]    reg_activation6_3_2;
wire[15:0]    reg_activation6_4_1;
wire[15:0]    reg_activation6_4_2;
wire[15:0]    reg_activation6_5_1;
wire[15:0]    reg_activation6_5_2;
wire[15:0]    reg_activation6_6_1;
wire[15:0]    reg_activation6_6_2;
wire[15:0]    reg_activation6_7_1;
wire[15:0]    reg_activation6_7_2;
wire[15:0]    reg_activation6_8_1;
wire[15:0]    reg_activation6_8_2;
wire[15:0]    reg_activation6_9_1;
wire[15:0]    reg_activation6_9_2;
wire[15:0]    reg_activation6_10_1;
wire[15:0]    reg_activation6_10_2;
wire[15:0]    reg_activation6_11_1;
wire[15:0]    reg_activation6_11_2;
wire[15:0]    reg_activation6_12_1;
wire[15:0]    reg_activation6_12_2;
wire[15:0]    reg_activation6_13_1;
wire[15:0]    reg_activation6_13_2;
wire[15:0]    reg_activation6_14_1;
wire[15:0]    reg_activation6_14_2;
wire[15:0]    reg_activation6_15_1;
wire[15:0]    reg_activation6_15_2;
wire[15:0]    reg_activation6_16_1;
wire[15:0]    reg_activation6_16_2;
wire[15:0]    reg_activation6_17_1;
wire[15:0]    reg_activation6_17_2;
wire[15:0]    reg_activation6_18_1;
wire[15:0]    reg_activation6_18_2;
wire[15:0]    reg_activation6_19_1;
wire[15:0]    reg_activation6_19_2;
wire[15:0]    reg_activation6_20_1;
wire[15:0]    reg_activation6_20_2;
wire[15:0]    reg_activation6_21_1;
wire[15:0]    reg_activation6_21_2;
wire[15:0]    reg_activation6_22_1;
wire[15:0]    reg_activation6_22_2;
wire[15:0]    reg_activation6_23_1;
wire[15:0]    reg_activation6_23_2;
wire[15:0]    reg_activation6_24_1;
wire[15:0]    reg_activation6_24_2;
wire[15:0]    reg_activation6_25_1;
wire[15:0]    reg_activation6_25_2;
wire[15:0]    reg_activation6_26_1;
wire[15:0]    reg_activation6_26_2;
wire[15:0]    reg_activation6_27_1;
wire[15:0]    reg_activation6_27_2;
wire[15:0]    reg_activation6_28_1;
wire[15:0]    reg_activation6_28_2;
wire[15:0]    reg_activation6_29_1;
wire[15:0]    reg_activation6_29_2;
wire[15:0]    reg_activation6_30_1;
wire[15:0]    reg_activation6_30_2;
wire[15:0]    reg_activation6_31_1;
wire[15:0]    reg_activation6_31_2;
wire[15:0]    reg_activation7_1_1;
wire[15:0]    reg_activation7_1_2;
wire[15:0]    reg_activation7_2_1;
wire[15:0]    reg_activation7_2_2;
wire[15:0]    reg_activation7_3_1;
wire[15:0]    reg_activation7_3_2;
wire[15:0]    reg_activation7_4_1;
wire[15:0]    reg_activation7_4_2;
wire[15:0]    reg_activation7_5_1;
wire[15:0]    reg_activation7_5_2;
wire[15:0]    reg_activation7_6_1;
wire[15:0]    reg_activation7_6_2;
wire[15:0]    reg_activation7_7_1;
wire[15:0]    reg_activation7_7_2;
wire[15:0]    reg_activation7_8_1;
wire[15:0]    reg_activation7_8_2;
wire[15:0]    reg_activation7_9_1;
wire[15:0]    reg_activation7_9_2;
wire[15:0]    reg_activation7_10_1;
wire[15:0]    reg_activation7_10_2;
wire[15:0]    reg_activation7_11_1;
wire[15:0]    reg_activation7_11_2;
wire[15:0]    reg_activation7_12_1;
wire[15:0]    reg_activation7_12_2;
wire[15:0]    reg_activation7_13_1;
wire[15:0]    reg_activation7_13_2;
wire[15:0]    reg_activation7_14_1;
wire[15:0]    reg_activation7_14_2;
wire[15:0]    reg_activation7_15_1;
wire[15:0]    reg_activation7_15_2;
wire[15:0]    reg_activation7_16_1;
wire[15:0]    reg_activation7_16_2;
wire[15:0]    reg_activation7_17_1;
wire[15:0]    reg_activation7_17_2;
wire[15:0]    reg_activation7_18_1;
wire[15:0]    reg_activation7_18_2;
wire[15:0]    reg_activation7_19_1;
wire[15:0]    reg_activation7_19_2;
wire[15:0]    reg_activation7_20_1;
wire[15:0]    reg_activation7_20_2;
wire[15:0]    reg_activation7_21_1;
wire[15:0]    reg_activation7_21_2;
wire[15:0]    reg_activation7_22_1;
wire[15:0]    reg_activation7_22_2;
wire[15:0]    reg_activation7_23_1;
wire[15:0]    reg_activation7_23_2;
wire[15:0]    reg_activation7_24_1;
wire[15:0]    reg_activation7_24_2;
wire[15:0]    reg_activation7_25_1;
wire[15:0]    reg_activation7_25_2;
wire[15:0]    reg_activation7_26_1;
wire[15:0]    reg_activation7_26_2;
wire[15:0]    reg_activation7_27_1;
wire[15:0]    reg_activation7_27_2;
wire[15:0]    reg_activation7_28_1;
wire[15:0]    reg_activation7_28_2;
wire[15:0]    reg_activation7_29_1;
wire[15:0]    reg_activation7_29_2;
wire[15:0]    reg_activation7_30_1;
wire[15:0]    reg_activation7_30_2;
wire[15:0]    reg_activation7_31_1;
wire[15:0]    reg_activation7_31_2;
wire[15:0]    reg_activation8_1_1;
wire[15:0]    reg_activation8_1_2;
wire[15:0]    reg_activation8_2_1;
wire[15:0]    reg_activation8_2_2;
wire[15:0]    reg_activation8_3_1;
wire[15:0]    reg_activation8_3_2;
wire[15:0]    reg_activation8_4_1;
wire[15:0]    reg_activation8_4_2;
wire[15:0]    reg_activation8_5_1;
wire[15:0]    reg_activation8_5_2;
wire[15:0]    reg_activation8_6_1;
wire[15:0]    reg_activation8_6_2;
wire[15:0]    reg_activation8_7_1;
wire[15:0]    reg_activation8_7_2;
wire[15:0]    reg_activation8_8_1;
wire[15:0]    reg_activation8_8_2;
wire[15:0]    reg_activation8_9_1;
wire[15:0]    reg_activation8_9_2;
wire[15:0]    reg_activation8_10_1;
wire[15:0]    reg_activation8_10_2;
wire[15:0]    reg_activation8_11_1;
wire[15:0]    reg_activation8_11_2;
wire[15:0]    reg_activation8_12_1;
wire[15:0]    reg_activation8_12_2;
wire[15:0]    reg_activation8_13_1;
wire[15:0]    reg_activation8_13_2;
wire[15:0]    reg_activation8_14_1;
wire[15:0]    reg_activation8_14_2;
wire[15:0]    reg_activation8_15_1;
wire[15:0]    reg_activation8_15_2;
wire[15:0]    reg_activation8_16_1;
wire[15:0]    reg_activation8_16_2;
wire[15:0]    reg_activation8_17_1;
wire[15:0]    reg_activation8_17_2;
wire[15:0]    reg_activation8_18_1;
wire[15:0]    reg_activation8_18_2;
wire[15:0]    reg_activation8_19_1;
wire[15:0]    reg_activation8_19_2;
wire[15:0]    reg_activation8_20_1;
wire[15:0]    reg_activation8_20_2;
wire[15:0]    reg_activation8_21_1;
wire[15:0]    reg_activation8_21_2;
wire[15:0]    reg_activation8_22_1;
wire[15:0]    reg_activation8_22_2;
wire[15:0]    reg_activation8_23_1;
wire[15:0]    reg_activation8_23_2;
wire[15:0]    reg_activation8_24_1;
wire[15:0]    reg_activation8_24_2;
wire[15:0]    reg_activation8_25_1;
wire[15:0]    reg_activation8_25_2;
wire[15:0]    reg_activation8_26_1;
wire[15:0]    reg_activation8_26_2;
wire[15:0]    reg_activation8_27_1;
wire[15:0]    reg_activation8_27_2;
wire[15:0]    reg_activation8_28_1;
wire[15:0]    reg_activation8_28_2;
wire[15:0]    reg_activation8_29_1;
wire[15:0]    reg_activation8_29_2;
wire[15:0]    reg_activation8_30_1;
wire[15:0]    reg_activation8_30_2;
wire[15:0]    reg_activation8_31_1;
wire[15:0]    reg_activation8_31_2;
wire[15:0]    reg_activation9_1_1;
wire[15:0]    reg_activation9_1_2;
wire[15:0]    reg_activation9_2_1;
wire[15:0]    reg_activation9_2_2;
wire[15:0]    reg_activation9_3_1;
wire[15:0]    reg_activation9_3_2;
wire[15:0]    reg_activation9_4_1;
wire[15:0]    reg_activation9_4_2;
wire[15:0]    reg_activation9_5_1;
wire[15:0]    reg_activation9_5_2;
wire[15:0]    reg_activation9_6_1;
wire[15:0]    reg_activation9_6_2;
wire[15:0]    reg_activation9_7_1;
wire[15:0]    reg_activation9_7_2;
wire[15:0]    reg_activation9_8_1;
wire[15:0]    reg_activation9_8_2;
wire[15:0]    reg_activation9_9_1;
wire[15:0]    reg_activation9_9_2;
wire[15:0]    reg_activation9_10_1;
wire[15:0]    reg_activation9_10_2;
wire[15:0]    reg_activation9_11_1;
wire[15:0]    reg_activation9_11_2;
wire[15:0]    reg_activation9_12_1;
wire[15:0]    reg_activation9_12_2;
wire[15:0]    reg_activation9_13_1;
wire[15:0]    reg_activation9_13_2;
wire[15:0]    reg_activation9_14_1;
wire[15:0]    reg_activation9_14_2;
wire[15:0]    reg_activation9_15_1;
wire[15:0]    reg_activation9_15_2;
wire[15:0]    reg_activation9_16_1;
wire[15:0]    reg_activation9_16_2;
wire[15:0]    reg_activation9_17_1;
wire[15:0]    reg_activation9_17_2;
wire[15:0]    reg_activation9_18_1;
wire[15:0]    reg_activation9_18_2;
wire[15:0]    reg_activation9_19_1;
wire[15:0]    reg_activation9_19_2;
wire[15:0]    reg_activation9_20_1;
wire[15:0]    reg_activation9_20_2;
wire[15:0]    reg_activation9_21_1;
wire[15:0]    reg_activation9_21_2;
wire[15:0]    reg_activation9_22_1;
wire[15:0]    reg_activation9_22_2;
wire[15:0]    reg_activation9_23_1;
wire[15:0]    reg_activation9_23_2;
wire[15:0]    reg_activation9_24_1;
wire[15:0]    reg_activation9_24_2;
wire[15:0]    reg_activation9_25_1;
wire[15:0]    reg_activation9_25_2;
wire[15:0]    reg_activation9_26_1;
wire[15:0]    reg_activation9_26_2;
wire[15:0]    reg_activation9_27_1;
wire[15:0]    reg_activation9_27_2;
wire[15:0]    reg_activation9_28_1;
wire[15:0]    reg_activation9_28_2;
wire[15:0]    reg_activation9_29_1;
wire[15:0]    reg_activation9_29_2;
wire[15:0]    reg_activation9_30_1;
wire[15:0]    reg_activation9_30_2;
wire[15:0]    reg_activation9_31_1;
wire[15:0]    reg_activation9_31_2;
wire[15:0]    reg_activation10_1_1;
wire[15:0]    reg_activation10_1_2;
wire[15:0]    reg_activation10_2_1;
wire[15:0]    reg_activation10_2_2;
wire[15:0]    reg_activation10_3_1;
wire[15:0]    reg_activation10_3_2;
wire[15:0]    reg_activation10_4_1;
wire[15:0]    reg_activation10_4_2;
wire[15:0]    reg_activation10_5_1;
wire[15:0]    reg_activation10_5_2;
wire[15:0]    reg_activation10_6_1;
wire[15:0]    reg_activation10_6_2;
wire[15:0]    reg_activation10_7_1;
wire[15:0]    reg_activation10_7_2;
wire[15:0]    reg_activation10_8_1;
wire[15:0]    reg_activation10_8_2;
wire[15:0]    reg_activation10_9_1;
wire[15:0]    reg_activation10_9_2;
wire[15:0]    reg_activation10_10_1;
wire[15:0]    reg_activation10_10_2;
wire[15:0]    reg_activation10_11_1;
wire[15:0]    reg_activation10_11_2;
wire[15:0]    reg_activation10_12_1;
wire[15:0]    reg_activation10_12_2;
wire[15:0]    reg_activation10_13_1;
wire[15:0]    reg_activation10_13_2;
wire[15:0]    reg_activation10_14_1;
wire[15:0]    reg_activation10_14_2;
wire[15:0]    reg_activation10_15_1;
wire[15:0]    reg_activation10_15_2;
wire[15:0]    reg_activation10_16_1;
wire[15:0]    reg_activation10_16_2;
wire[15:0]    reg_activation10_17_1;
wire[15:0]    reg_activation10_17_2;
wire[15:0]    reg_activation10_18_1;
wire[15:0]    reg_activation10_18_2;
wire[15:0]    reg_activation10_19_1;
wire[15:0]    reg_activation10_19_2;
wire[15:0]    reg_activation10_20_1;
wire[15:0]    reg_activation10_20_2;
wire[15:0]    reg_activation10_21_1;
wire[15:0]    reg_activation10_21_2;
wire[15:0]    reg_activation10_22_1;
wire[15:0]    reg_activation10_22_2;
wire[15:0]    reg_activation10_23_1;
wire[15:0]    reg_activation10_23_2;
wire[15:0]    reg_activation10_24_1;
wire[15:0]    reg_activation10_24_2;
wire[15:0]    reg_activation10_25_1;
wire[15:0]    reg_activation10_25_2;
wire[15:0]    reg_activation10_26_1;
wire[15:0]    reg_activation10_26_2;
wire[15:0]    reg_activation10_27_1;
wire[15:0]    reg_activation10_27_2;
wire[15:0]    reg_activation10_28_1;
wire[15:0]    reg_activation10_28_2;
wire[15:0]    reg_activation10_29_1;
wire[15:0]    reg_activation10_29_2;
wire[15:0]    reg_activation10_30_1;
wire[15:0]    reg_activation10_30_2;
wire[15:0]    reg_activation10_31_1;
wire[15:0]    reg_activation10_31_2;
wire[15:0]    reg_activation11_1_1;
wire[15:0]    reg_activation11_1_2;
wire[15:0]    reg_activation11_2_1;
wire[15:0]    reg_activation11_2_2;
wire[15:0]    reg_activation11_3_1;
wire[15:0]    reg_activation11_3_2;
wire[15:0]    reg_activation11_4_1;
wire[15:0]    reg_activation11_4_2;
wire[15:0]    reg_activation11_5_1;
wire[15:0]    reg_activation11_5_2;
wire[15:0]    reg_activation11_6_1;
wire[15:0]    reg_activation11_6_2;
wire[15:0]    reg_activation11_7_1;
wire[15:0]    reg_activation11_7_2;
wire[15:0]    reg_activation11_8_1;
wire[15:0]    reg_activation11_8_2;
wire[15:0]    reg_activation11_9_1;
wire[15:0]    reg_activation11_9_2;
wire[15:0]    reg_activation11_10_1;
wire[15:0]    reg_activation11_10_2;
wire[15:0]    reg_activation11_11_1;
wire[15:0]    reg_activation11_11_2;
wire[15:0]    reg_activation11_12_1;
wire[15:0]    reg_activation11_12_2;
wire[15:0]    reg_activation11_13_1;
wire[15:0]    reg_activation11_13_2;
wire[15:0]    reg_activation11_14_1;
wire[15:0]    reg_activation11_14_2;
wire[15:0]    reg_activation11_15_1;
wire[15:0]    reg_activation11_15_2;
wire[15:0]    reg_activation11_16_1;
wire[15:0]    reg_activation11_16_2;
wire[15:0]    reg_activation11_17_1;
wire[15:0]    reg_activation11_17_2;
wire[15:0]    reg_activation11_18_1;
wire[15:0]    reg_activation11_18_2;
wire[15:0]    reg_activation11_19_1;
wire[15:0]    reg_activation11_19_2;
wire[15:0]    reg_activation11_20_1;
wire[15:0]    reg_activation11_20_2;
wire[15:0]    reg_activation11_21_1;
wire[15:0]    reg_activation11_21_2;
wire[15:0]    reg_activation11_22_1;
wire[15:0]    reg_activation11_22_2;
wire[15:0]    reg_activation11_23_1;
wire[15:0]    reg_activation11_23_2;
wire[15:0]    reg_activation11_24_1;
wire[15:0]    reg_activation11_24_2;
wire[15:0]    reg_activation11_25_1;
wire[15:0]    reg_activation11_25_2;
wire[15:0]    reg_activation11_26_1;
wire[15:0]    reg_activation11_26_2;
wire[15:0]    reg_activation11_27_1;
wire[15:0]    reg_activation11_27_2;
wire[15:0]    reg_activation11_28_1;
wire[15:0]    reg_activation11_28_2;
wire[15:0]    reg_activation11_29_1;
wire[15:0]    reg_activation11_29_2;
wire[15:0]    reg_activation11_30_1;
wire[15:0]    reg_activation11_30_2;
wire[15:0]    reg_activation11_31_1;
wire[15:0]    reg_activation11_31_2;
wire[15:0]    reg_activation12_1_1;
wire[15:0]    reg_activation12_1_2;
wire[15:0]    reg_activation12_2_1;
wire[15:0]    reg_activation12_2_2;
wire[15:0]    reg_activation12_3_1;
wire[15:0]    reg_activation12_3_2;
wire[15:0]    reg_activation12_4_1;
wire[15:0]    reg_activation12_4_2;
wire[15:0]    reg_activation12_5_1;
wire[15:0]    reg_activation12_5_2;
wire[15:0]    reg_activation12_6_1;
wire[15:0]    reg_activation12_6_2;
wire[15:0]    reg_activation12_7_1;
wire[15:0]    reg_activation12_7_2;
wire[15:0]    reg_activation12_8_1;
wire[15:0]    reg_activation12_8_2;
wire[15:0]    reg_activation12_9_1;
wire[15:0]    reg_activation12_9_2;
wire[15:0]    reg_activation12_10_1;
wire[15:0]    reg_activation12_10_2;
wire[15:0]    reg_activation12_11_1;
wire[15:0]    reg_activation12_11_2;
wire[15:0]    reg_activation12_12_1;
wire[15:0]    reg_activation12_12_2;
wire[15:0]    reg_activation12_13_1;
wire[15:0]    reg_activation12_13_2;
wire[15:0]    reg_activation12_14_1;
wire[15:0]    reg_activation12_14_2;
wire[15:0]    reg_activation12_15_1;
wire[15:0]    reg_activation12_15_2;
wire[15:0]    reg_activation12_16_1;
wire[15:0]    reg_activation12_16_2;
wire[15:0]    reg_activation12_17_1;
wire[15:0]    reg_activation12_17_2;
wire[15:0]    reg_activation12_18_1;
wire[15:0]    reg_activation12_18_2;
wire[15:0]    reg_activation12_19_1;
wire[15:0]    reg_activation12_19_2;
wire[15:0]    reg_activation12_20_1;
wire[15:0]    reg_activation12_20_2;
wire[15:0]    reg_activation12_21_1;
wire[15:0]    reg_activation12_21_2;
wire[15:0]    reg_activation12_22_1;
wire[15:0]    reg_activation12_22_2;
wire[15:0]    reg_activation12_23_1;
wire[15:0]    reg_activation12_23_2;
wire[15:0]    reg_activation12_24_1;
wire[15:0]    reg_activation12_24_2;
wire[15:0]    reg_activation12_25_1;
wire[15:0]    reg_activation12_25_2;
wire[15:0]    reg_activation12_26_1;
wire[15:0]    reg_activation12_26_2;
wire[15:0]    reg_activation12_27_1;
wire[15:0]    reg_activation12_27_2;
wire[15:0]    reg_activation12_28_1;
wire[15:0]    reg_activation12_28_2;
wire[15:0]    reg_activation12_29_1;
wire[15:0]    reg_activation12_29_2;
wire[15:0]    reg_activation12_30_1;
wire[15:0]    reg_activation12_30_2;
wire[15:0]    reg_activation12_31_1;
wire[15:0]    reg_activation12_31_2;
wire[15:0]    reg_activation13_1_1;
wire[15:0]    reg_activation13_1_2;
wire[15:0]    reg_activation13_2_1;
wire[15:0]    reg_activation13_2_2;
wire[15:0]    reg_activation13_3_1;
wire[15:0]    reg_activation13_3_2;
wire[15:0]    reg_activation13_4_1;
wire[15:0]    reg_activation13_4_2;
wire[15:0]    reg_activation13_5_1;
wire[15:0]    reg_activation13_5_2;
wire[15:0]    reg_activation13_6_1;
wire[15:0]    reg_activation13_6_2;
wire[15:0]    reg_activation13_7_1;
wire[15:0]    reg_activation13_7_2;
wire[15:0]    reg_activation13_8_1;
wire[15:0]    reg_activation13_8_2;
wire[15:0]    reg_activation13_9_1;
wire[15:0]    reg_activation13_9_2;
wire[15:0]    reg_activation13_10_1;
wire[15:0]    reg_activation13_10_2;
wire[15:0]    reg_activation13_11_1;
wire[15:0]    reg_activation13_11_2;
wire[15:0]    reg_activation13_12_1;
wire[15:0]    reg_activation13_12_2;
wire[15:0]    reg_activation13_13_1;
wire[15:0]    reg_activation13_13_2;
wire[15:0]    reg_activation13_14_1;
wire[15:0]    reg_activation13_14_2;
wire[15:0]    reg_activation13_15_1;
wire[15:0]    reg_activation13_15_2;
wire[15:0]    reg_activation13_16_1;
wire[15:0]    reg_activation13_16_2;
wire[15:0]    reg_activation13_17_1;
wire[15:0]    reg_activation13_17_2;
wire[15:0]    reg_activation13_18_1;
wire[15:0]    reg_activation13_18_2;
wire[15:0]    reg_activation13_19_1;
wire[15:0]    reg_activation13_19_2;
wire[15:0]    reg_activation13_20_1;
wire[15:0]    reg_activation13_20_2;
wire[15:0]    reg_activation13_21_1;
wire[15:0]    reg_activation13_21_2;
wire[15:0]    reg_activation13_22_1;
wire[15:0]    reg_activation13_22_2;
wire[15:0]    reg_activation13_23_1;
wire[15:0]    reg_activation13_23_2;
wire[15:0]    reg_activation13_24_1;
wire[15:0]    reg_activation13_24_2;
wire[15:0]    reg_activation13_25_1;
wire[15:0]    reg_activation13_25_2;
wire[15:0]    reg_activation13_26_1;
wire[15:0]    reg_activation13_26_2;
wire[15:0]    reg_activation13_27_1;
wire[15:0]    reg_activation13_27_2;
wire[15:0]    reg_activation13_28_1;
wire[15:0]    reg_activation13_28_2;
wire[15:0]    reg_activation13_29_1;
wire[15:0]    reg_activation13_29_2;
wire[15:0]    reg_activation13_30_1;
wire[15:0]    reg_activation13_30_2;
wire[15:0]    reg_activation13_31_1;
wire[15:0]    reg_activation13_31_2;
wire[15:0]    reg_activation14_1_1;
wire[15:0]    reg_activation14_1_2;
wire[15:0]    reg_activation14_2_1;
wire[15:0]    reg_activation14_2_2;
wire[15:0]    reg_activation14_3_1;
wire[15:0]    reg_activation14_3_2;
wire[15:0]    reg_activation14_4_1;
wire[15:0]    reg_activation14_4_2;
wire[15:0]    reg_activation14_5_1;
wire[15:0]    reg_activation14_5_2;
wire[15:0]    reg_activation14_6_1;
wire[15:0]    reg_activation14_6_2;
wire[15:0]    reg_activation14_7_1;
wire[15:0]    reg_activation14_7_2;
wire[15:0]    reg_activation14_8_1;
wire[15:0]    reg_activation14_8_2;
wire[15:0]    reg_activation14_9_1;
wire[15:0]    reg_activation14_9_2;
wire[15:0]    reg_activation14_10_1;
wire[15:0]    reg_activation14_10_2;
wire[15:0]    reg_activation14_11_1;
wire[15:0]    reg_activation14_11_2;
wire[15:0]    reg_activation14_12_1;
wire[15:0]    reg_activation14_12_2;
wire[15:0]    reg_activation14_13_1;
wire[15:0]    reg_activation14_13_2;
wire[15:0]    reg_activation14_14_1;
wire[15:0]    reg_activation14_14_2;
wire[15:0]    reg_activation14_15_1;
wire[15:0]    reg_activation14_15_2;
wire[15:0]    reg_activation14_16_1;
wire[15:0]    reg_activation14_16_2;
wire[15:0]    reg_activation14_17_1;
wire[15:0]    reg_activation14_17_2;
wire[15:0]    reg_activation14_18_1;
wire[15:0]    reg_activation14_18_2;
wire[15:0]    reg_activation14_19_1;
wire[15:0]    reg_activation14_19_2;
wire[15:0]    reg_activation14_20_1;
wire[15:0]    reg_activation14_20_2;
wire[15:0]    reg_activation14_21_1;
wire[15:0]    reg_activation14_21_2;
wire[15:0]    reg_activation14_22_1;
wire[15:0]    reg_activation14_22_2;
wire[15:0]    reg_activation14_23_1;
wire[15:0]    reg_activation14_23_2;
wire[15:0]    reg_activation14_24_1;
wire[15:0]    reg_activation14_24_2;
wire[15:0]    reg_activation14_25_1;
wire[15:0]    reg_activation14_25_2;
wire[15:0]    reg_activation14_26_1;
wire[15:0]    reg_activation14_26_2;
wire[15:0]    reg_activation14_27_1;
wire[15:0]    reg_activation14_27_2;
wire[15:0]    reg_activation14_28_1;
wire[15:0]    reg_activation14_28_2;
wire[15:0]    reg_activation14_29_1;
wire[15:0]    reg_activation14_29_2;
wire[15:0]    reg_activation14_30_1;
wire[15:0]    reg_activation14_30_2;
wire[15:0]    reg_activation14_31_1;
wire[15:0]    reg_activation14_31_2;
wire[15:0]    reg_activation15_1_1;
wire[15:0]    reg_activation15_1_2;
wire[15:0]    reg_activation15_2_1;
wire[15:0]    reg_activation15_2_2;
wire[15:0]    reg_activation15_3_1;
wire[15:0]    reg_activation15_3_2;
wire[15:0]    reg_activation15_4_1;
wire[15:0]    reg_activation15_4_2;
wire[15:0]    reg_activation15_5_1;
wire[15:0]    reg_activation15_5_2;
wire[15:0]    reg_activation15_6_1;
wire[15:0]    reg_activation15_6_2;
wire[15:0]    reg_activation15_7_1;
wire[15:0]    reg_activation15_7_2;
wire[15:0]    reg_activation15_8_1;
wire[15:0]    reg_activation15_8_2;
wire[15:0]    reg_activation15_9_1;
wire[15:0]    reg_activation15_9_2;
wire[15:0]    reg_activation15_10_1;
wire[15:0]    reg_activation15_10_2;
wire[15:0]    reg_activation15_11_1;
wire[15:0]    reg_activation15_11_2;
wire[15:0]    reg_activation15_12_1;
wire[15:0]    reg_activation15_12_2;
wire[15:0]    reg_activation15_13_1;
wire[15:0]    reg_activation15_13_2;
wire[15:0]    reg_activation15_14_1;
wire[15:0]    reg_activation15_14_2;
wire[15:0]    reg_activation15_15_1;
wire[15:0]    reg_activation15_15_2;
wire[15:0]    reg_activation15_16_1;
wire[15:0]    reg_activation15_16_2;
wire[15:0]    reg_activation15_17_1;
wire[15:0]    reg_activation15_17_2;
wire[15:0]    reg_activation15_18_1;
wire[15:0]    reg_activation15_18_2;
wire[15:0]    reg_activation15_19_1;
wire[15:0]    reg_activation15_19_2;
wire[15:0]    reg_activation15_20_1;
wire[15:0]    reg_activation15_20_2;
wire[15:0]    reg_activation15_21_1;
wire[15:0]    reg_activation15_21_2;
wire[15:0]    reg_activation15_22_1;
wire[15:0]    reg_activation15_22_2;
wire[15:0]    reg_activation15_23_1;
wire[15:0]    reg_activation15_23_2;
wire[15:0]    reg_activation15_24_1;
wire[15:0]    reg_activation15_24_2;
wire[15:0]    reg_activation15_25_1;
wire[15:0]    reg_activation15_25_2;
wire[15:0]    reg_activation15_26_1;
wire[15:0]    reg_activation15_26_2;
wire[15:0]    reg_activation15_27_1;
wire[15:0]    reg_activation15_27_2;
wire[15:0]    reg_activation15_28_1;
wire[15:0]    reg_activation15_28_2;
wire[15:0]    reg_activation15_29_1;
wire[15:0]    reg_activation15_29_2;
wire[15:0]    reg_activation15_30_1;
wire[15:0]    reg_activation15_30_2;
wire[15:0]    reg_activation15_31_1;
wire[15:0]    reg_activation15_31_2;
wire[15:0]    reg_activation16_1_1;
wire[15:0]    reg_activation16_1_2;
wire[15:0]    reg_activation16_2_1;
wire[15:0]    reg_activation16_2_2;
wire[15:0]    reg_activation16_3_1;
wire[15:0]    reg_activation16_3_2;
wire[15:0]    reg_activation16_4_1;
wire[15:0]    reg_activation16_4_2;
wire[15:0]    reg_activation16_5_1;
wire[15:0]    reg_activation16_5_2;
wire[15:0]    reg_activation16_6_1;
wire[15:0]    reg_activation16_6_2;
wire[15:0]    reg_activation16_7_1;
wire[15:0]    reg_activation16_7_2;
wire[15:0]    reg_activation16_8_1;
wire[15:0]    reg_activation16_8_2;
wire[15:0]    reg_activation16_9_1;
wire[15:0]    reg_activation16_9_2;
wire[15:0]    reg_activation16_10_1;
wire[15:0]    reg_activation16_10_2;
wire[15:0]    reg_activation16_11_1;
wire[15:0]    reg_activation16_11_2;
wire[15:0]    reg_activation16_12_1;
wire[15:0]    reg_activation16_12_2;
wire[15:0]    reg_activation16_13_1;
wire[15:0]    reg_activation16_13_2;
wire[15:0]    reg_activation16_14_1;
wire[15:0]    reg_activation16_14_2;
wire[15:0]    reg_activation16_15_1;
wire[15:0]    reg_activation16_15_2;
wire[15:0]    reg_activation16_16_1;
wire[15:0]    reg_activation16_16_2;
wire[15:0]    reg_activation16_17_1;
wire[15:0]    reg_activation16_17_2;
wire[15:0]    reg_activation16_18_1;
wire[15:0]    reg_activation16_18_2;
wire[15:0]    reg_activation16_19_1;
wire[15:0]    reg_activation16_19_2;
wire[15:0]    reg_activation16_20_1;
wire[15:0]    reg_activation16_20_2;
wire[15:0]    reg_activation16_21_1;
wire[15:0]    reg_activation16_21_2;
wire[15:0]    reg_activation16_22_1;
wire[15:0]    reg_activation16_22_2;
wire[15:0]    reg_activation16_23_1;
wire[15:0]    reg_activation16_23_2;
wire[15:0]    reg_activation16_24_1;
wire[15:0]    reg_activation16_24_2;
wire[15:0]    reg_activation16_25_1;
wire[15:0]    reg_activation16_25_2;
wire[15:0]    reg_activation16_26_1;
wire[15:0]    reg_activation16_26_2;
wire[15:0]    reg_activation16_27_1;
wire[15:0]    reg_activation16_27_2;
wire[15:0]    reg_activation16_28_1;
wire[15:0]    reg_activation16_28_2;
wire[15:0]    reg_activation16_29_1;
wire[15:0]    reg_activation16_29_2;
wire[15:0]    reg_activation16_30_1;
wire[15:0]    reg_activation16_30_2;
wire[15:0]    reg_activation16_31_1;
wire[15:0]    reg_activation16_31_2;
wire[15:0]    reg_activation17_1_1;
wire[15:0]    reg_activation17_1_2;
wire[15:0]    reg_activation17_2_1;
wire[15:0]    reg_activation17_2_2;
wire[15:0]    reg_activation17_3_1;
wire[15:0]    reg_activation17_3_2;
wire[15:0]    reg_activation17_4_1;
wire[15:0]    reg_activation17_4_2;
wire[15:0]    reg_activation17_5_1;
wire[15:0]    reg_activation17_5_2;
wire[15:0]    reg_activation17_6_1;
wire[15:0]    reg_activation17_6_2;
wire[15:0]    reg_activation17_7_1;
wire[15:0]    reg_activation17_7_2;
wire[15:0]    reg_activation17_8_1;
wire[15:0]    reg_activation17_8_2;
wire[15:0]    reg_activation17_9_1;
wire[15:0]    reg_activation17_9_2;
wire[15:0]    reg_activation17_10_1;
wire[15:0]    reg_activation17_10_2;
wire[15:0]    reg_activation17_11_1;
wire[15:0]    reg_activation17_11_2;
wire[15:0]    reg_activation17_12_1;
wire[15:0]    reg_activation17_12_2;
wire[15:0]    reg_activation17_13_1;
wire[15:0]    reg_activation17_13_2;
wire[15:0]    reg_activation17_14_1;
wire[15:0]    reg_activation17_14_2;
wire[15:0]    reg_activation17_15_1;
wire[15:0]    reg_activation17_15_2;
wire[15:0]    reg_activation17_16_1;
wire[15:0]    reg_activation17_16_2;
wire[15:0]    reg_activation17_17_1;
wire[15:0]    reg_activation17_17_2;
wire[15:0]    reg_activation17_18_1;
wire[15:0]    reg_activation17_18_2;
wire[15:0]    reg_activation17_19_1;
wire[15:0]    reg_activation17_19_2;
wire[15:0]    reg_activation17_20_1;
wire[15:0]    reg_activation17_20_2;
wire[15:0]    reg_activation17_21_1;
wire[15:0]    reg_activation17_21_2;
wire[15:0]    reg_activation17_22_1;
wire[15:0]    reg_activation17_22_2;
wire[15:0]    reg_activation17_23_1;
wire[15:0]    reg_activation17_23_2;
wire[15:0]    reg_activation17_24_1;
wire[15:0]    reg_activation17_24_2;
wire[15:0]    reg_activation17_25_1;
wire[15:0]    reg_activation17_25_2;
wire[15:0]    reg_activation17_26_1;
wire[15:0]    reg_activation17_26_2;
wire[15:0]    reg_activation17_27_1;
wire[15:0]    reg_activation17_27_2;
wire[15:0]    reg_activation17_28_1;
wire[15:0]    reg_activation17_28_2;
wire[15:0]    reg_activation17_29_1;
wire[15:0]    reg_activation17_29_2;
wire[15:0]    reg_activation17_30_1;
wire[15:0]    reg_activation17_30_2;
wire[15:0]    reg_activation17_31_1;
wire[15:0]    reg_activation17_31_2;
wire[15:0]    reg_activation18_1_1;
wire[15:0]    reg_activation18_1_2;
wire[15:0]    reg_activation18_2_1;
wire[15:0]    reg_activation18_2_2;
wire[15:0]    reg_activation18_3_1;
wire[15:0]    reg_activation18_3_2;
wire[15:0]    reg_activation18_4_1;
wire[15:0]    reg_activation18_4_2;
wire[15:0]    reg_activation18_5_1;
wire[15:0]    reg_activation18_5_2;
wire[15:0]    reg_activation18_6_1;
wire[15:0]    reg_activation18_6_2;
wire[15:0]    reg_activation18_7_1;
wire[15:0]    reg_activation18_7_2;
wire[15:0]    reg_activation18_8_1;
wire[15:0]    reg_activation18_8_2;
wire[15:0]    reg_activation18_9_1;
wire[15:0]    reg_activation18_9_2;
wire[15:0]    reg_activation18_10_1;
wire[15:0]    reg_activation18_10_2;
wire[15:0]    reg_activation18_11_1;
wire[15:0]    reg_activation18_11_2;
wire[15:0]    reg_activation18_12_1;
wire[15:0]    reg_activation18_12_2;
wire[15:0]    reg_activation18_13_1;
wire[15:0]    reg_activation18_13_2;
wire[15:0]    reg_activation18_14_1;
wire[15:0]    reg_activation18_14_2;
wire[15:0]    reg_activation18_15_1;
wire[15:0]    reg_activation18_15_2;
wire[15:0]    reg_activation18_16_1;
wire[15:0]    reg_activation18_16_2;
wire[15:0]    reg_activation18_17_1;
wire[15:0]    reg_activation18_17_2;
wire[15:0]    reg_activation18_18_1;
wire[15:0]    reg_activation18_18_2;
wire[15:0]    reg_activation18_19_1;
wire[15:0]    reg_activation18_19_2;
wire[15:0]    reg_activation18_20_1;
wire[15:0]    reg_activation18_20_2;
wire[15:0]    reg_activation18_21_1;
wire[15:0]    reg_activation18_21_2;
wire[15:0]    reg_activation18_22_1;
wire[15:0]    reg_activation18_22_2;
wire[15:0]    reg_activation18_23_1;
wire[15:0]    reg_activation18_23_2;
wire[15:0]    reg_activation18_24_1;
wire[15:0]    reg_activation18_24_2;
wire[15:0]    reg_activation18_25_1;
wire[15:0]    reg_activation18_25_2;
wire[15:0]    reg_activation18_26_1;
wire[15:0]    reg_activation18_26_2;
wire[15:0]    reg_activation18_27_1;
wire[15:0]    reg_activation18_27_2;
wire[15:0]    reg_activation18_28_1;
wire[15:0]    reg_activation18_28_2;
wire[15:0]    reg_activation18_29_1;
wire[15:0]    reg_activation18_29_2;
wire[15:0]    reg_activation18_30_1;
wire[15:0]    reg_activation18_30_2;
wire[15:0]    reg_activation18_31_1;
wire[15:0]    reg_activation18_31_2;
wire[15:0]    reg_activation19_1_1;
wire[15:0]    reg_activation19_1_2;
wire[15:0]    reg_activation19_2_1;
wire[15:0]    reg_activation19_2_2;
wire[15:0]    reg_activation19_3_1;
wire[15:0]    reg_activation19_3_2;
wire[15:0]    reg_activation19_4_1;
wire[15:0]    reg_activation19_4_2;
wire[15:0]    reg_activation19_5_1;
wire[15:0]    reg_activation19_5_2;
wire[15:0]    reg_activation19_6_1;
wire[15:0]    reg_activation19_6_2;
wire[15:0]    reg_activation19_7_1;
wire[15:0]    reg_activation19_7_2;
wire[15:0]    reg_activation19_8_1;
wire[15:0]    reg_activation19_8_2;
wire[15:0]    reg_activation19_9_1;
wire[15:0]    reg_activation19_9_2;
wire[15:0]    reg_activation19_10_1;
wire[15:0]    reg_activation19_10_2;
wire[15:0]    reg_activation19_11_1;
wire[15:0]    reg_activation19_11_2;
wire[15:0]    reg_activation19_12_1;
wire[15:0]    reg_activation19_12_2;
wire[15:0]    reg_activation19_13_1;
wire[15:0]    reg_activation19_13_2;
wire[15:0]    reg_activation19_14_1;
wire[15:0]    reg_activation19_14_2;
wire[15:0]    reg_activation19_15_1;
wire[15:0]    reg_activation19_15_2;
wire[15:0]    reg_activation19_16_1;
wire[15:0]    reg_activation19_16_2;
wire[15:0]    reg_activation19_17_1;
wire[15:0]    reg_activation19_17_2;
wire[15:0]    reg_activation19_18_1;
wire[15:0]    reg_activation19_18_2;
wire[15:0]    reg_activation19_19_1;
wire[15:0]    reg_activation19_19_2;
wire[15:0]    reg_activation19_20_1;
wire[15:0]    reg_activation19_20_2;
wire[15:0]    reg_activation19_21_1;
wire[15:0]    reg_activation19_21_2;
wire[15:0]    reg_activation19_22_1;
wire[15:0]    reg_activation19_22_2;
wire[15:0]    reg_activation19_23_1;
wire[15:0]    reg_activation19_23_2;
wire[15:0]    reg_activation19_24_1;
wire[15:0]    reg_activation19_24_2;
wire[15:0]    reg_activation19_25_1;
wire[15:0]    reg_activation19_25_2;
wire[15:0]    reg_activation19_26_1;
wire[15:0]    reg_activation19_26_2;
wire[15:0]    reg_activation19_27_1;
wire[15:0]    reg_activation19_27_2;
wire[15:0]    reg_activation19_28_1;
wire[15:0]    reg_activation19_28_2;
wire[15:0]    reg_activation19_29_1;
wire[15:0]    reg_activation19_29_2;
wire[15:0]    reg_activation19_30_1;
wire[15:0]    reg_activation19_30_2;
wire[15:0]    reg_activation19_31_1;
wire[15:0]    reg_activation19_31_2;
wire[15:0]    reg_activation20_1_1;
wire[15:0]    reg_activation20_1_2;
wire[15:0]    reg_activation20_2_1;
wire[15:0]    reg_activation20_2_2;
wire[15:0]    reg_activation20_3_1;
wire[15:0]    reg_activation20_3_2;
wire[15:0]    reg_activation20_4_1;
wire[15:0]    reg_activation20_4_2;
wire[15:0]    reg_activation20_5_1;
wire[15:0]    reg_activation20_5_2;
wire[15:0]    reg_activation20_6_1;
wire[15:0]    reg_activation20_6_2;
wire[15:0]    reg_activation20_7_1;
wire[15:0]    reg_activation20_7_2;
wire[15:0]    reg_activation20_8_1;
wire[15:0]    reg_activation20_8_2;
wire[15:0]    reg_activation20_9_1;
wire[15:0]    reg_activation20_9_2;
wire[15:0]    reg_activation20_10_1;
wire[15:0]    reg_activation20_10_2;
wire[15:0]    reg_activation20_11_1;
wire[15:0]    reg_activation20_11_2;
wire[15:0]    reg_activation20_12_1;
wire[15:0]    reg_activation20_12_2;
wire[15:0]    reg_activation20_13_1;
wire[15:0]    reg_activation20_13_2;
wire[15:0]    reg_activation20_14_1;
wire[15:0]    reg_activation20_14_2;
wire[15:0]    reg_activation20_15_1;
wire[15:0]    reg_activation20_15_2;
wire[15:0]    reg_activation20_16_1;
wire[15:0]    reg_activation20_16_2;
wire[15:0]    reg_activation20_17_1;
wire[15:0]    reg_activation20_17_2;
wire[15:0]    reg_activation20_18_1;
wire[15:0]    reg_activation20_18_2;
wire[15:0]    reg_activation20_19_1;
wire[15:0]    reg_activation20_19_2;
wire[15:0]    reg_activation20_20_1;
wire[15:0]    reg_activation20_20_2;
wire[15:0]    reg_activation20_21_1;
wire[15:0]    reg_activation20_21_2;
wire[15:0]    reg_activation20_22_1;
wire[15:0]    reg_activation20_22_2;
wire[15:0]    reg_activation20_23_1;
wire[15:0]    reg_activation20_23_2;
wire[15:0]    reg_activation20_24_1;
wire[15:0]    reg_activation20_24_2;
wire[15:0]    reg_activation20_25_1;
wire[15:0]    reg_activation20_25_2;
wire[15:0]    reg_activation20_26_1;
wire[15:0]    reg_activation20_26_2;
wire[15:0]    reg_activation20_27_1;
wire[15:0]    reg_activation20_27_2;
wire[15:0]    reg_activation20_28_1;
wire[15:0]    reg_activation20_28_2;
wire[15:0]    reg_activation20_29_1;
wire[15:0]    reg_activation20_29_2;
wire[15:0]    reg_activation20_30_1;
wire[15:0]    reg_activation20_30_2;
wire[15:0]    reg_activation20_31_1;
wire[15:0]    reg_activation20_31_2;
wire[15:0]    reg_activation21_1_1;
wire[15:0]    reg_activation21_1_2;
wire[15:0]    reg_activation21_2_1;
wire[15:0]    reg_activation21_2_2;
wire[15:0]    reg_activation21_3_1;
wire[15:0]    reg_activation21_3_2;
wire[15:0]    reg_activation21_4_1;
wire[15:0]    reg_activation21_4_2;
wire[15:0]    reg_activation21_5_1;
wire[15:0]    reg_activation21_5_2;
wire[15:0]    reg_activation21_6_1;
wire[15:0]    reg_activation21_6_2;
wire[15:0]    reg_activation21_7_1;
wire[15:0]    reg_activation21_7_2;
wire[15:0]    reg_activation21_8_1;
wire[15:0]    reg_activation21_8_2;
wire[15:0]    reg_activation21_9_1;
wire[15:0]    reg_activation21_9_2;
wire[15:0]    reg_activation21_10_1;
wire[15:0]    reg_activation21_10_2;
wire[15:0]    reg_activation21_11_1;
wire[15:0]    reg_activation21_11_2;
wire[15:0]    reg_activation21_12_1;
wire[15:0]    reg_activation21_12_2;
wire[15:0]    reg_activation21_13_1;
wire[15:0]    reg_activation21_13_2;
wire[15:0]    reg_activation21_14_1;
wire[15:0]    reg_activation21_14_2;
wire[15:0]    reg_activation21_15_1;
wire[15:0]    reg_activation21_15_2;
wire[15:0]    reg_activation21_16_1;
wire[15:0]    reg_activation21_16_2;
wire[15:0]    reg_activation21_17_1;
wire[15:0]    reg_activation21_17_2;
wire[15:0]    reg_activation21_18_1;
wire[15:0]    reg_activation21_18_2;
wire[15:0]    reg_activation21_19_1;
wire[15:0]    reg_activation21_19_2;
wire[15:0]    reg_activation21_20_1;
wire[15:0]    reg_activation21_20_2;
wire[15:0]    reg_activation21_21_1;
wire[15:0]    reg_activation21_21_2;
wire[15:0]    reg_activation21_22_1;
wire[15:0]    reg_activation21_22_2;
wire[15:0]    reg_activation21_23_1;
wire[15:0]    reg_activation21_23_2;
wire[15:0]    reg_activation21_24_1;
wire[15:0]    reg_activation21_24_2;
wire[15:0]    reg_activation21_25_1;
wire[15:0]    reg_activation21_25_2;
wire[15:0]    reg_activation21_26_1;
wire[15:0]    reg_activation21_26_2;
wire[15:0]    reg_activation21_27_1;
wire[15:0]    reg_activation21_27_2;
wire[15:0]    reg_activation21_28_1;
wire[15:0]    reg_activation21_28_2;
wire[15:0]    reg_activation21_29_1;
wire[15:0]    reg_activation21_29_2;
wire[15:0]    reg_activation21_30_1;
wire[15:0]    reg_activation21_30_2;
wire[15:0]    reg_activation21_31_1;
wire[15:0]    reg_activation21_31_2;
wire[15:0]    reg_activation22_1_1;
wire[15:0]    reg_activation22_1_2;
wire[15:0]    reg_activation22_2_1;
wire[15:0]    reg_activation22_2_2;
wire[15:0]    reg_activation22_3_1;
wire[15:0]    reg_activation22_3_2;
wire[15:0]    reg_activation22_4_1;
wire[15:0]    reg_activation22_4_2;
wire[15:0]    reg_activation22_5_1;
wire[15:0]    reg_activation22_5_2;
wire[15:0]    reg_activation22_6_1;
wire[15:0]    reg_activation22_6_2;
wire[15:0]    reg_activation22_7_1;
wire[15:0]    reg_activation22_7_2;
wire[15:0]    reg_activation22_8_1;
wire[15:0]    reg_activation22_8_2;
wire[15:0]    reg_activation22_9_1;
wire[15:0]    reg_activation22_9_2;
wire[15:0]    reg_activation22_10_1;
wire[15:0]    reg_activation22_10_2;
wire[15:0]    reg_activation22_11_1;
wire[15:0]    reg_activation22_11_2;
wire[15:0]    reg_activation22_12_1;
wire[15:0]    reg_activation22_12_2;
wire[15:0]    reg_activation22_13_1;
wire[15:0]    reg_activation22_13_2;
wire[15:0]    reg_activation22_14_1;
wire[15:0]    reg_activation22_14_2;
wire[15:0]    reg_activation22_15_1;
wire[15:0]    reg_activation22_15_2;
wire[15:0]    reg_activation22_16_1;
wire[15:0]    reg_activation22_16_2;
wire[15:0]    reg_activation22_17_1;
wire[15:0]    reg_activation22_17_2;
wire[15:0]    reg_activation22_18_1;
wire[15:0]    reg_activation22_18_2;
wire[15:0]    reg_activation22_19_1;
wire[15:0]    reg_activation22_19_2;
wire[15:0]    reg_activation22_20_1;
wire[15:0]    reg_activation22_20_2;
wire[15:0]    reg_activation22_21_1;
wire[15:0]    reg_activation22_21_2;
wire[15:0]    reg_activation22_22_1;
wire[15:0]    reg_activation22_22_2;
wire[15:0]    reg_activation22_23_1;
wire[15:0]    reg_activation22_23_2;
wire[15:0]    reg_activation22_24_1;
wire[15:0]    reg_activation22_24_2;
wire[15:0]    reg_activation22_25_1;
wire[15:0]    reg_activation22_25_2;
wire[15:0]    reg_activation22_26_1;
wire[15:0]    reg_activation22_26_2;
wire[15:0]    reg_activation22_27_1;
wire[15:0]    reg_activation22_27_2;
wire[15:0]    reg_activation22_28_1;
wire[15:0]    reg_activation22_28_2;
wire[15:0]    reg_activation22_29_1;
wire[15:0]    reg_activation22_29_2;
wire[15:0]    reg_activation22_30_1;
wire[15:0]    reg_activation22_30_2;
wire[15:0]    reg_activation22_31_1;
wire[15:0]    reg_activation22_31_2;
wire[15:0]    reg_activation23_1_1;
wire[15:0]    reg_activation23_1_2;
wire[15:0]    reg_activation23_2_1;
wire[15:0]    reg_activation23_2_2;
wire[15:0]    reg_activation23_3_1;
wire[15:0]    reg_activation23_3_2;
wire[15:0]    reg_activation23_4_1;
wire[15:0]    reg_activation23_4_2;
wire[15:0]    reg_activation23_5_1;
wire[15:0]    reg_activation23_5_2;
wire[15:0]    reg_activation23_6_1;
wire[15:0]    reg_activation23_6_2;
wire[15:0]    reg_activation23_7_1;
wire[15:0]    reg_activation23_7_2;
wire[15:0]    reg_activation23_8_1;
wire[15:0]    reg_activation23_8_2;
wire[15:0]    reg_activation23_9_1;
wire[15:0]    reg_activation23_9_2;
wire[15:0]    reg_activation23_10_1;
wire[15:0]    reg_activation23_10_2;
wire[15:0]    reg_activation23_11_1;
wire[15:0]    reg_activation23_11_2;
wire[15:0]    reg_activation23_12_1;
wire[15:0]    reg_activation23_12_2;
wire[15:0]    reg_activation23_13_1;
wire[15:0]    reg_activation23_13_2;
wire[15:0]    reg_activation23_14_1;
wire[15:0]    reg_activation23_14_2;
wire[15:0]    reg_activation23_15_1;
wire[15:0]    reg_activation23_15_2;
wire[15:0]    reg_activation23_16_1;
wire[15:0]    reg_activation23_16_2;
wire[15:0]    reg_activation23_17_1;
wire[15:0]    reg_activation23_17_2;
wire[15:0]    reg_activation23_18_1;
wire[15:0]    reg_activation23_18_2;
wire[15:0]    reg_activation23_19_1;
wire[15:0]    reg_activation23_19_2;
wire[15:0]    reg_activation23_20_1;
wire[15:0]    reg_activation23_20_2;
wire[15:0]    reg_activation23_21_1;
wire[15:0]    reg_activation23_21_2;
wire[15:0]    reg_activation23_22_1;
wire[15:0]    reg_activation23_22_2;
wire[15:0]    reg_activation23_23_1;
wire[15:0]    reg_activation23_23_2;
wire[15:0]    reg_activation23_24_1;
wire[15:0]    reg_activation23_24_2;
wire[15:0]    reg_activation23_25_1;
wire[15:0]    reg_activation23_25_2;
wire[15:0]    reg_activation23_26_1;
wire[15:0]    reg_activation23_26_2;
wire[15:0]    reg_activation23_27_1;
wire[15:0]    reg_activation23_27_2;
wire[15:0]    reg_activation23_28_1;
wire[15:0]    reg_activation23_28_2;
wire[15:0]    reg_activation23_29_1;
wire[15:0]    reg_activation23_29_2;
wire[15:0]    reg_activation23_30_1;
wire[15:0]    reg_activation23_30_2;
wire[15:0]    reg_activation23_31_1;
wire[15:0]    reg_activation23_31_2;
wire[15:0]    reg_activation24_1_1;
wire[15:0]    reg_activation24_1_2;
wire[15:0]    reg_activation24_2_1;
wire[15:0]    reg_activation24_2_2;
wire[15:0]    reg_activation24_3_1;
wire[15:0]    reg_activation24_3_2;
wire[15:0]    reg_activation24_4_1;
wire[15:0]    reg_activation24_4_2;
wire[15:0]    reg_activation24_5_1;
wire[15:0]    reg_activation24_5_2;
wire[15:0]    reg_activation24_6_1;
wire[15:0]    reg_activation24_6_2;
wire[15:0]    reg_activation24_7_1;
wire[15:0]    reg_activation24_7_2;
wire[15:0]    reg_activation24_8_1;
wire[15:0]    reg_activation24_8_2;
wire[15:0]    reg_activation24_9_1;
wire[15:0]    reg_activation24_9_2;
wire[15:0]    reg_activation24_10_1;
wire[15:0]    reg_activation24_10_2;
wire[15:0]    reg_activation24_11_1;
wire[15:0]    reg_activation24_11_2;
wire[15:0]    reg_activation24_12_1;
wire[15:0]    reg_activation24_12_2;
wire[15:0]    reg_activation24_13_1;
wire[15:0]    reg_activation24_13_2;
wire[15:0]    reg_activation24_14_1;
wire[15:0]    reg_activation24_14_2;
wire[15:0]    reg_activation24_15_1;
wire[15:0]    reg_activation24_15_2;
wire[15:0]    reg_activation24_16_1;
wire[15:0]    reg_activation24_16_2;
wire[15:0]    reg_activation24_17_1;
wire[15:0]    reg_activation24_17_2;
wire[15:0]    reg_activation24_18_1;
wire[15:0]    reg_activation24_18_2;
wire[15:0]    reg_activation24_19_1;
wire[15:0]    reg_activation24_19_2;
wire[15:0]    reg_activation24_20_1;
wire[15:0]    reg_activation24_20_2;
wire[15:0]    reg_activation24_21_1;
wire[15:0]    reg_activation24_21_2;
wire[15:0]    reg_activation24_22_1;
wire[15:0]    reg_activation24_22_2;
wire[15:0]    reg_activation24_23_1;
wire[15:0]    reg_activation24_23_2;
wire[15:0]    reg_activation24_24_1;
wire[15:0]    reg_activation24_24_2;
wire[15:0]    reg_activation24_25_1;
wire[15:0]    reg_activation24_25_2;
wire[15:0]    reg_activation24_26_1;
wire[15:0]    reg_activation24_26_2;
wire[15:0]    reg_activation24_27_1;
wire[15:0]    reg_activation24_27_2;
wire[15:0]    reg_activation24_28_1;
wire[15:0]    reg_activation24_28_2;
wire[15:0]    reg_activation24_29_1;
wire[15:0]    reg_activation24_29_2;
wire[15:0]    reg_activation24_30_1;
wire[15:0]    reg_activation24_30_2;
wire[15:0]    reg_activation24_31_1;
wire[15:0]    reg_activation24_31_2;
wire[15:0]    reg_activation25_1_1;
wire[15:0]    reg_activation25_1_2;
wire[15:0]    reg_activation25_2_1;
wire[15:0]    reg_activation25_2_2;
wire[15:0]    reg_activation25_3_1;
wire[15:0]    reg_activation25_3_2;
wire[15:0]    reg_activation25_4_1;
wire[15:0]    reg_activation25_4_2;
wire[15:0]    reg_activation25_5_1;
wire[15:0]    reg_activation25_5_2;
wire[15:0]    reg_activation25_6_1;
wire[15:0]    reg_activation25_6_2;
wire[15:0]    reg_activation25_7_1;
wire[15:0]    reg_activation25_7_2;
wire[15:0]    reg_activation25_8_1;
wire[15:0]    reg_activation25_8_2;
wire[15:0]    reg_activation25_9_1;
wire[15:0]    reg_activation25_9_2;
wire[15:0]    reg_activation25_10_1;
wire[15:0]    reg_activation25_10_2;
wire[15:0]    reg_activation25_11_1;
wire[15:0]    reg_activation25_11_2;
wire[15:0]    reg_activation25_12_1;
wire[15:0]    reg_activation25_12_2;
wire[15:0]    reg_activation25_13_1;
wire[15:0]    reg_activation25_13_2;
wire[15:0]    reg_activation25_14_1;
wire[15:0]    reg_activation25_14_2;
wire[15:0]    reg_activation25_15_1;
wire[15:0]    reg_activation25_15_2;
wire[15:0]    reg_activation25_16_1;
wire[15:0]    reg_activation25_16_2;
wire[15:0]    reg_activation25_17_1;
wire[15:0]    reg_activation25_17_2;
wire[15:0]    reg_activation25_18_1;
wire[15:0]    reg_activation25_18_2;
wire[15:0]    reg_activation25_19_1;
wire[15:0]    reg_activation25_19_2;
wire[15:0]    reg_activation25_20_1;
wire[15:0]    reg_activation25_20_2;
wire[15:0]    reg_activation25_21_1;
wire[15:0]    reg_activation25_21_2;
wire[15:0]    reg_activation25_22_1;
wire[15:0]    reg_activation25_22_2;
wire[15:0]    reg_activation25_23_1;
wire[15:0]    reg_activation25_23_2;
wire[15:0]    reg_activation25_24_1;
wire[15:0]    reg_activation25_24_2;
wire[15:0]    reg_activation25_25_1;
wire[15:0]    reg_activation25_25_2;
wire[15:0]    reg_activation25_26_1;
wire[15:0]    reg_activation25_26_2;
wire[15:0]    reg_activation25_27_1;
wire[15:0]    reg_activation25_27_2;
wire[15:0]    reg_activation25_28_1;
wire[15:0]    reg_activation25_28_2;
wire[15:0]    reg_activation25_29_1;
wire[15:0]    reg_activation25_29_2;
wire[15:0]    reg_activation25_30_1;
wire[15:0]    reg_activation25_30_2;
wire[15:0]    reg_activation25_31_1;
wire[15:0]    reg_activation25_31_2;
wire[15:0]    reg_activation26_1_1;
wire[15:0]    reg_activation26_1_2;
wire[15:0]    reg_activation26_2_1;
wire[15:0]    reg_activation26_2_2;
wire[15:0]    reg_activation26_3_1;
wire[15:0]    reg_activation26_3_2;
wire[15:0]    reg_activation26_4_1;
wire[15:0]    reg_activation26_4_2;
wire[15:0]    reg_activation26_5_1;
wire[15:0]    reg_activation26_5_2;
wire[15:0]    reg_activation26_6_1;
wire[15:0]    reg_activation26_6_2;
wire[15:0]    reg_activation26_7_1;
wire[15:0]    reg_activation26_7_2;
wire[15:0]    reg_activation26_8_1;
wire[15:0]    reg_activation26_8_2;
wire[15:0]    reg_activation26_9_1;
wire[15:0]    reg_activation26_9_2;
wire[15:0]    reg_activation26_10_1;
wire[15:0]    reg_activation26_10_2;
wire[15:0]    reg_activation26_11_1;
wire[15:0]    reg_activation26_11_2;
wire[15:0]    reg_activation26_12_1;
wire[15:0]    reg_activation26_12_2;
wire[15:0]    reg_activation26_13_1;
wire[15:0]    reg_activation26_13_2;
wire[15:0]    reg_activation26_14_1;
wire[15:0]    reg_activation26_14_2;
wire[15:0]    reg_activation26_15_1;
wire[15:0]    reg_activation26_15_2;
wire[15:0]    reg_activation26_16_1;
wire[15:0]    reg_activation26_16_2;
wire[15:0]    reg_activation26_17_1;
wire[15:0]    reg_activation26_17_2;
wire[15:0]    reg_activation26_18_1;
wire[15:0]    reg_activation26_18_2;
wire[15:0]    reg_activation26_19_1;
wire[15:0]    reg_activation26_19_2;
wire[15:0]    reg_activation26_20_1;
wire[15:0]    reg_activation26_20_2;
wire[15:0]    reg_activation26_21_1;
wire[15:0]    reg_activation26_21_2;
wire[15:0]    reg_activation26_22_1;
wire[15:0]    reg_activation26_22_2;
wire[15:0]    reg_activation26_23_1;
wire[15:0]    reg_activation26_23_2;
wire[15:0]    reg_activation26_24_1;
wire[15:0]    reg_activation26_24_2;
wire[15:0]    reg_activation26_25_1;
wire[15:0]    reg_activation26_25_2;
wire[15:0]    reg_activation26_26_1;
wire[15:0]    reg_activation26_26_2;
wire[15:0]    reg_activation26_27_1;
wire[15:0]    reg_activation26_27_2;
wire[15:0]    reg_activation26_28_1;
wire[15:0]    reg_activation26_28_2;
wire[15:0]    reg_activation26_29_1;
wire[15:0]    reg_activation26_29_2;
wire[15:0]    reg_activation26_30_1;
wire[15:0]    reg_activation26_30_2;
wire[15:0]    reg_activation26_31_1;
wire[15:0]    reg_activation26_31_2;
wire[15:0]    reg_activation27_1_1;
wire[15:0]    reg_activation27_1_2;
wire[15:0]    reg_activation27_2_1;
wire[15:0]    reg_activation27_2_2;
wire[15:0]    reg_activation27_3_1;
wire[15:0]    reg_activation27_3_2;
wire[15:0]    reg_activation27_4_1;
wire[15:0]    reg_activation27_4_2;
wire[15:0]    reg_activation27_5_1;
wire[15:0]    reg_activation27_5_2;
wire[15:0]    reg_activation27_6_1;
wire[15:0]    reg_activation27_6_2;
wire[15:0]    reg_activation27_7_1;
wire[15:0]    reg_activation27_7_2;
wire[15:0]    reg_activation27_8_1;
wire[15:0]    reg_activation27_8_2;
wire[15:0]    reg_activation27_9_1;
wire[15:0]    reg_activation27_9_2;
wire[15:0]    reg_activation27_10_1;
wire[15:0]    reg_activation27_10_2;
wire[15:0]    reg_activation27_11_1;
wire[15:0]    reg_activation27_11_2;
wire[15:0]    reg_activation27_12_1;
wire[15:0]    reg_activation27_12_2;
wire[15:0]    reg_activation27_13_1;
wire[15:0]    reg_activation27_13_2;
wire[15:0]    reg_activation27_14_1;
wire[15:0]    reg_activation27_14_2;
wire[15:0]    reg_activation27_15_1;
wire[15:0]    reg_activation27_15_2;
wire[15:0]    reg_activation27_16_1;
wire[15:0]    reg_activation27_16_2;
wire[15:0]    reg_activation27_17_1;
wire[15:0]    reg_activation27_17_2;
wire[15:0]    reg_activation27_18_1;
wire[15:0]    reg_activation27_18_2;
wire[15:0]    reg_activation27_19_1;
wire[15:0]    reg_activation27_19_2;
wire[15:0]    reg_activation27_20_1;
wire[15:0]    reg_activation27_20_2;
wire[15:0]    reg_activation27_21_1;
wire[15:0]    reg_activation27_21_2;
wire[15:0]    reg_activation27_22_1;
wire[15:0]    reg_activation27_22_2;
wire[15:0]    reg_activation27_23_1;
wire[15:0]    reg_activation27_23_2;
wire[15:0]    reg_activation27_24_1;
wire[15:0]    reg_activation27_24_2;
wire[15:0]    reg_activation27_25_1;
wire[15:0]    reg_activation27_25_2;
wire[15:0]    reg_activation27_26_1;
wire[15:0]    reg_activation27_26_2;
wire[15:0]    reg_activation27_27_1;
wire[15:0]    reg_activation27_27_2;
wire[15:0]    reg_activation27_28_1;
wire[15:0]    reg_activation27_28_2;
wire[15:0]    reg_activation27_29_1;
wire[15:0]    reg_activation27_29_2;
wire[15:0]    reg_activation27_30_1;
wire[15:0]    reg_activation27_30_2;
wire[15:0]    reg_activation27_31_1;
wire[15:0]    reg_activation27_31_2;
wire[15:0]    reg_activation28_1_1;
wire[15:0]    reg_activation28_1_2;
wire[15:0]    reg_activation28_2_1;
wire[15:0]    reg_activation28_2_2;
wire[15:0]    reg_activation28_3_1;
wire[15:0]    reg_activation28_3_2;
wire[15:0]    reg_activation28_4_1;
wire[15:0]    reg_activation28_4_2;
wire[15:0]    reg_activation28_5_1;
wire[15:0]    reg_activation28_5_2;
wire[15:0]    reg_activation28_6_1;
wire[15:0]    reg_activation28_6_2;
wire[15:0]    reg_activation28_7_1;
wire[15:0]    reg_activation28_7_2;
wire[15:0]    reg_activation28_8_1;
wire[15:0]    reg_activation28_8_2;
wire[15:0]    reg_activation28_9_1;
wire[15:0]    reg_activation28_9_2;
wire[15:0]    reg_activation28_10_1;
wire[15:0]    reg_activation28_10_2;
wire[15:0]    reg_activation28_11_1;
wire[15:0]    reg_activation28_11_2;
wire[15:0]    reg_activation28_12_1;
wire[15:0]    reg_activation28_12_2;
wire[15:0]    reg_activation28_13_1;
wire[15:0]    reg_activation28_13_2;
wire[15:0]    reg_activation28_14_1;
wire[15:0]    reg_activation28_14_2;
wire[15:0]    reg_activation28_15_1;
wire[15:0]    reg_activation28_15_2;
wire[15:0]    reg_activation28_16_1;
wire[15:0]    reg_activation28_16_2;
wire[15:0]    reg_activation28_17_1;
wire[15:0]    reg_activation28_17_2;
wire[15:0]    reg_activation28_18_1;
wire[15:0]    reg_activation28_18_2;
wire[15:0]    reg_activation28_19_1;
wire[15:0]    reg_activation28_19_2;
wire[15:0]    reg_activation28_20_1;
wire[15:0]    reg_activation28_20_2;
wire[15:0]    reg_activation28_21_1;
wire[15:0]    reg_activation28_21_2;
wire[15:0]    reg_activation28_22_1;
wire[15:0]    reg_activation28_22_2;
wire[15:0]    reg_activation28_23_1;
wire[15:0]    reg_activation28_23_2;
wire[15:0]    reg_activation28_24_1;
wire[15:0]    reg_activation28_24_2;
wire[15:0]    reg_activation28_25_1;
wire[15:0]    reg_activation28_25_2;
wire[15:0]    reg_activation28_26_1;
wire[15:0]    reg_activation28_26_2;
wire[15:0]    reg_activation28_27_1;
wire[15:0]    reg_activation28_27_2;
wire[15:0]    reg_activation28_28_1;
wire[15:0]    reg_activation28_28_2;
wire[15:0]    reg_activation28_29_1;
wire[15:0]    reg_activation28_29_2;
wire[15:0]    reg_activation28_30_1;
wire[15:0]    reg_activation28_30_2;
wire[15:0]    reg_activation28_31_1;
wire[15:0]    reg_activation28_31_2;
wire[15:0]    reg_activation29_1_1;
wire[15:0]    reg_activation29_1_2;
wire[15:0]    reg_activation29_2_1;
wire[15:0]    reg_activation29_2_2;
wire[15:0]    reg_activation29_3_1;
wire[15:0]    reg_activation29_3_2;
wire[15:0]    reg_activation29_4_1;
wire[15:0]    reg_activation29_4_2;
wire[15:0]    reg_activation29_5_1;
wire[15:0]    reg_activation29_5_2;
wire[15:0]    reg_activation29_6_1;
wire[15:0]    reg_activation29_6_2;
wire[15:0]    reg_activation29_7_1;
wire[15:0]    reg_activation29_7_2;
wire[15:0]    reg_activation29_8_1;
wire[15:0]    reg_activation29_8_2;
wire[15:0]    reg_activation29_9_1;
wire[15:0]    reg_activation29_9_2;
wire[15:0]    reg_activation29_10_1;
wire[15:0]    reg_activation29_10_2;
wire[15:0]    reg_activation29_11_1;
wire[15:0]    reg_activation29_11_2;
wire[15:0]    reg_activation29_12_1;
wire[15:0]    reg_activation29_12_2;
wire[15:0]    reg_activation29_13_1;
wire[15:0]    reg_activation29_13_2;
wire[15:0]    reg_activation29_14_1;
wire[15:0]    reg_activation29_14_2;
wire[15:0]    reg_activation29_15_1;
wire[15:0]    reg_activation29_15_2;
wire[15:0]    reg_activation29_16_1;
wire[15:0]    reg_activation29_16_2;
wire[15:0]    reg_activation29_17_1;
wire[15:0]    reg_activation29_17_2;
wire[15:0]    reg_activation29_18_1;
wire[15:0]    reg_activation29_18_2;
wire[15:0]    reg_activation29_19_1;
wire[15:0]    reg_activation29_19_2;
wire[15:0]    reg_activation29_20_1;
wire[15:0]    reg_activation29_20_2;
wire[15:0]    reg_activation29_21_1;
wire[15:0]    reg_activation29_21_2;
wire[15:0]    reg_activation29_22_1;
wire[15:0]    reg_activation29_22_2;
wire[15:0]    reg_activation29_23_1;
wire[15:0]    reg_activation29_23_2;
wire[15:0]    reg_activation29_24_1;
wire[15:0]    reg_activation29_24_2;
wire[15:0]    reg_activation29_25_1;
wire[15:0]    reg_activation29_25_2;
wire[15:0]    reg_activation29_26_1;
wire[15:0]    reg_activation29_26_2;
wire[15:0]    reg_activation29_27_1;
wire[15:0]    reg_activation29_27_2;
wire[15:0]    reg_activation29_28_1;
wire[15:0]    reg_activation29_28_2;
wire[15:0]    reg_activation29_29_1;
wire[15:0]    reg_activation29_29_2;
wire[15:0]    reg_activation29_30_1;
wire[15:0]    reg_activation29_30_2;
wire[15:0]    reg_activation29_31_1;
wire[15:0]    reg_activation29_31_2;
wire[15:0]    reg_activation30_1_1;
wire[15:0]    reg_activation30_1_2;
wire[15:0]    reg_activation30_2_1;
wire[15:0]    reg_activation30_2_2;
wire[15:0]    reg_activation30_3_1;
wire[15:0]    reg_activation30_3_2;
wire[15:0]    reg_activation30_4_1;
wire[15:0]    reg_activation30_4_2;
wire[15:0]    reg_activation30_5_1;
wire[15:0]    reg_activation30_5_2;
wire[15:0]    reg_activation30_6_1;
wire[15:0]    reg_activation30_6_2;
wire[15:0]    reg_activation30_7_1;
wire[15:0]    reg_activation30_7_2;
wire[15:0]    reg_activation30_8_1;
wire[15:0]    reg_activation30_8_2;
wire[15:0]    reg_activation30_9_1;
wire[15:0]    reg_activation30_9_2;
wire[15:0]    reg_activation30_10_1;
wire[15:0]    reg_activation30_10_2;
wire[15:0]    reg_activation30_11_1;
wire[15:0]    reg_activation30_11_2;
wire[15:0]    reg_activation30_12_1;
wire[15:0]    reg_activation30_12_2;
wire[15:0]    reg_activation30_13_1;
wire[15:0]    reg_activation30_13_2;
wire[15:0]    reg_activation30_14_1;
wire[15:0]    reg_activation30_14_2;
wire[15:0]    reg_activation30_15_1;
wire[15:0]    reg_activation30_15_2;
wire[15:0]    reg_activation30_16_1;
wire[15:0]    reg_activation30_16_2;
wire[15:0]    reg_activation30_17_1;
wire[15:0]    reg_activation30_17_2;
wire[15:0]    reg_activation30_18_1;
wire[15:0]    reg_activation30_18_2;
wire[15:0]    reg_activation30_19_1;
wire[15:0]    reg_activation30_19_2;
wire[15:0]    reg_activation30_20_1;
wire[15:0]    reg_activation30_20_2;
wire[15:0]    reg_activation30_21_1;
wire[15:0]    reg_activation30_21_2;
wire[15:0]    reg_activation30_22_1;
wire[15:0]    reg_activation30_22_2;
wire[15:0]    reg_activation30_23_1;
wire[15:0]    reg_activation30_23_2;
wire[15:0]    reg_activation30_24_1;
wire[15:0]    reg_activation30_24_2;
wire[15:0]    reg_activation30_25_1;
wire[15:0]    reg_activation30_25_2;
wire[15:0]    reg_activation30_26_1;
wire[15:0]    reg_activation30_26_2;
wire[15:0]    reg_activation30_27_1;
wire[15:0]    reg_activation30_27_2;
wire[15:0]    reg_activation30_28_1;
wire[15:0]    reg_activation30_28_2;
wire[15:0]    reg_activation30_29_1;
wire[15:0]    reg_activation30_29_2;
wire[15:0]    reg_activation30_30_1;
wire[15:0]    reg_activation30_30_2;
wire[15:0]    reg_activation30_31_1;
wire[15:0]    reg_activation30_31_2;
wire[15:0]    reg_activation31_1_1;
wire[15:0]    reg_activation31_1_2;
wire[15:0]    reg_activation31_2_1;
wire[15:0]    reg_activation31_2_2;
wire[15:0]    reg_activation31_3_1;
wire[15:0]    reg_activation31_3_2;
wire[15:0]    reg_activation31_4_1;
wire[15:0]    reg_activation31_4_2;
wire[15:0]    reg_activation31_5_1;
wire[15:0]    reg_activation31_5_2;
wire[15:0]    reg_activation31_6_1;
wire[15:0]    reg_activation31_6_2;
wire[15:0]    reg_activation31_7_1;
wire[15:0]    reg_activation31_7_2;
wire[15:0]    reg_activation31_8_1;
wire[15:0]    reg_activation31_8_2;
wire[15:0]    reg_activation31_9_1;
wire[15:0]    reg_activation31_9_2;
wire[15:0]    reg_activation31_10_1;
wire[15:0]    reg_activation31_10_2;
wire[15:0]    reg_activation31_11_1;
wire[15:0]    reg_activation31_11_2;
wire[15:0]    reg_activation31_12_1;
wire[15:0]    reg_activation31_12_2;
wire[15:0]    reg_activation31_13_1;
wire[15:0]    reg_activation31_13_2;
wire[15:0]    reg_activation31_14_1;
wire[15:0]    reg_activation31_14_2;
wire[15:0]    reg_activation31_15_1;
wire[15:0]    reg_activation31_15_2;
wire[15:0]    reg_activation31_16_1;
wire[15:0]    reg_activation31_16_2;
wire[15:0]    reg_activation31_17_1;
wire[15:0]    reg_activation31_17_2;
wire[15:0]    reg_activation31_18_1;
wire[15:0]    reg_activation31_18_2;
wire[15:0]    reg_activation31_19_1;
wire[15:0]    reg_activation31_19_2;
wire[15:0]    reg_activation31_20_1;
wire[15:0]    reg_activation31_20_2;
wire[15:0]    reg_activation31_21_1;
wire[15:0]    reg_activation31_21_2;
wire[15:0]    reg_activation31_22_1;
wire[15:0]    reg_activation31_22_2;
wire[15:0]    reg_activation31_23_1;
wire[15:0]    reg_activation31_23_2;
wire[15:0]    reg_activation31_24_1;
wire[15:0]    reg_activation31_24_2;
wire[15:0]    reg_activation31_25_1;
wire[15:0]    reg_activation31_25_2;
wire[15:0]    reg_activation31_26_1;
wire[15:0]    reg_activation31_26_2;
wire[15:0]    reg_activation31_27_1;
wire[15:0]    reg_activation31_27_2;
wire[15:0]    reg_activation31_28_1;
wire[15:0]    reg_activation31_28_2;
wire[15:0]    reg_activation31_29_1;
wire[15:0]    reg_activation31_29_2;
wire[15:0]    reg_activation31_30_1;
wire[15:0]    reg_activation31_30_2;
wire[15:0]    reg_activation31_31_1;
wire[15:0]    reg_activation31_31_2;
wire[15:0]    reg_activation32_1_1;
wire[15:0]    reg_activation32_1_2;
wire[15:0]    reg_activation32_2_1;
wire[15:0]    reg_activation32_2_2;
wire[15:0]    reg_activation32_3_1;
wire[15:0]    reg_activation32_3_2;
wire[15:0]    reg_activation32_4_1;
wire[15:0]    reg_activation32_4_2;
wire[15:0]    reg_activation32_5_1;
wire[15:0]    reg_activation32_5_2;
wire[15:0]    reg_activation32_6_1;
wire[15:0]    reg_activation32_6_2;
wire[15:0]    reg_activation32_7_1;
wire[15:0]    reg_activation32_7_2;
wire[15:0]    reg_activation32_8_1;
wire[15:0]    reg_activation32_8_2;
wire[15:0]    reg_activation32_9_1;
wire[15:0]    reg_activation32_9_2;
wire[15:0]    reg_activation32_10_1;
wire[15:0]    reg_activation32_10_2;
wire[15:0]    reg_activation32_11_1;
wire[15:0]    reg_activation32_11_2;
wire[15:0]    reg_activation32_12_1;
wire[15:0]    reg_activation32_12_2;
wire[15:0]    reg_activation32_13_1;
wire[15:0]    reg_activation32_13_2;
wire[15:0]    reg_activation32_14_1;
wire[15:0]    reg_activation32_14_2;
wire[15:0]    reg_activation32_15_1;
wire[15:0]    reg_activation32_15_2;
wire[15:0]    reg_activation32_16_1;
wire[15:0]    reg_activation32_16_2;
wire[15:0]    reg_activation32_17_1;
wire[15:0]    reg_activation32_17_2;
wire[15:0]    reg_activation32_18_1;
wire[15:0]    reg_activation32_18_2;
wire[15:0]    reg_activation32_19_1;
wire[15:0]    reg_activation32_19_2;
wire[15:0]    reg_activation32_20_1;
wire[15:0]    reg_activation32_20_2;
wire[15:0]    reg_activation32_21_1;
wire[15:0]    reg_activation32_21_2;
wire[15:0]    reg_activation32_22_1;
wire[15:0]    reg_activation32_22_2;
wire[15:0]    reg_activation32_23_1;
wire[15:0]    reg_activation32_23_2;
wire[15:0]    reg_activation32_24_1;
wire[15:0]    reg_activation32_24_2;
wire[15:0]    reg_activation32_25_1;
wire[15:0]    reg_activation32_25_2;
wire[15:0]    reg_activation32_26_1;
wire[15:0]    reg_activation32_26_2;
wire[15:0]    reg_activation32_27_1;
wire[15:0]    reg_activation32_27_2;
wire[15:0]    reg_activation32_28_1;
wire[15:0]    reg_activation32_28_2;
wire[15:0]    reg_activation32_29_1;
wire[15:0]    reg_activation32_29_2;
wire[15:0]    reg_activation32_30_1;
wire[15:0]    reg_activation32_30_2;
wire[15:0]    reg_activation32_31_1;
wire[15:0]    reg_activation32_31_2;
wire[15:0]    reg_weight1_1_1;
wire[15:0]    reg_psum1_1_1;
wire[15:0]    reg_weight1_1_2;
wire[15:0]    reg_psum1_1_2;
wire[15:0]    reg_weight1_2_1;
wire[15:0]    reg_psum1_2_1;
wire[15:0]    reg_weight1_2_2;
wire[15:0]    reg_psum1_2_2;
wire[15:0]    reg_weight1_3_1;
wire[15:0]    reg_psum1_3_1;
wire[15:0]    reg_weight1_3_2;
wire[15:0]    reg_psum1_3_2;
wire[15:0]    reg_weight1_4_1;
wire[15:0]    reg_psum1_4_1;
wire[15:0]    reg_weight1_4_2;
wire[15:0]    reg_psum1_4_2;
wire[15:0]    reg_weight1_5_1;
wire[15:0]    reg_psum1_5_1;
wire[15:0]    reg_weight1_5_2;
wire[15:0]    reg_psum1_5_2;
wire[15:0]    reg_weight1_6_1;
wire[15:0]    reg_psum1_6_1;
wire[15:0]    reg_weight1_6_2;
wire[15:0]    reg_psum1_6_2;
wire[15:0]    reg_weight1_7_1;
wire[15:0]    reg_psum1_7_1;
wire[15:0]    reg_weight1_7_2;
wire[15:0]    reg_psum1_7_2;
wire[15:0]    reg_weight1_8_1;
wire[15:0]    reg_psum1_8_1;
wire[15:0]    reg_weight1_8_2;
wire[15:0]    reg_psum1_8_2;
wire[15:0]    reg_weight1_9_1;
wire[15:0]    reg_psum1_9_1;
wire[15:0]    reg_weight1_9_2;
wire[15:0]    reg_psum1_9_2;
wire[15:0]    reg_weight1_10_1;
wire[15:0]    reg_psum1_10_1;
wire[15:0]    reg_weight1_10_2;
wire[15:0]    reg_psum1_10_2;
wire[15:0]    reg_weight1_11_1;
wire[15:0]    reg_psum1_11_1;
wire[15:0]    reg_weight1_11_2;
wire[15:0]    reg_psum1_11_2;
wire[15:0]    reg_weight1_12_1;
wire[15:0]    reg_psum1_12_1;
wire[15:0]    reg_weight1_12_2;
wire[15:0]    reg_psum1_12_2;
wire[15:0]    reg_weight1_13_1;
wire[15:0]    reg_psum1_13_1;
wire[15:0]    reg_weight1_13_2;
wire[15:0]    reg_psum1_13_2;
wire[15:0]    reg_weight1_14_1;
wire[15:0]    reg_psum1_14_1;
wire[15:0]    reg_weight1_14_2;
wire[15:0]    reg_psum1_14_2;
wire[15:0]    reg_weight1_15_1;
wire[15:0]    reg_psum1_15_1;
wire[15:0]    reg_weight1_15_2;
wire[15:0]    reg_psum1_15_2;
wire[15:0]    reg_weight1_16_1;
wire[15:0]    reg_psum1_16_1;
wire[15:0]    reg_weight1_16_2;
wire[15:0]    reg_psum1_16_2;
wire[15:0]    reg_weight1_17_1;
wire[15:0]    reg_psum1_17_1;
wire[15:0]    reg_weight1_17_2;
wire[15:0]    reg_psum1_17_2;
wire[15:0]    reg_weight1_18_1;
wire[15:0]    reg_psum1_18_1;
wire[15:0]    reg_weight1_18_2;
wire[15:0]    reg_psum1_18_2;
wire[15:0]    reg_weight1_19_1;
wire[15:0]    reg_psum1_19_1;
wire[15:0]    reg_weight1_19_2;
wire[15:0]    reg_psum1_19_2;
wire[15:0]    reg_weight1_20_1;
wire[15:0]    reg_psum1_20_1;
wire[15:0]    reg_weight1_20_2;
wire[15:0]    reg_psum1_20_2;
wire[15:0]    reg_weight1_21_1;
wire[15:0]    reg_psum1_21_1;
wire[15:0]    reg_weight1_21_2;
wire[15:0]    reg_psum1_21_2;
wire[15:0]    reg_weight1_22_1;
wire[15:0]    reg_psum1_22_1;
wire[15:0]    reg_weight1_22_2;
wire[15:0]    reg_psum1_22_2;
wire[15:0]    reg_weight1_23_1;
wire[15:0]    reg_psum1_23_1;
wire[15:0]    reg_weight1_23_2;
wire[15:0]    reg_psum1_23_2;
wire[15:0]    reg_weight1_24_1;
wire[15:0]    reg_psum1_24_1;
wire[15:0]    reg_weight1_24_2;
wire[15:0]    reg_psum1_24_2;
wire[15:0]    reg_weight1_25_1;
wire[15:0]    reg_psum1_25_1;
wire[15:0]    reg_weight1_25_2;
wire[15:0]    reg_psum1_25_2;
wire[15:0]    reg_weight1_26_1;
wire[15:0]    reg_psum1_26_1;
wire[15:0]    reg_weight1_26_2;
wire[15:0]    reg_psum1_26_2;
wire[15:0]    reg_weight1_27_1;
wire[15:0]    reg_psum1_27_1;
wire[15:0]    reg_weight1_27_2;
wire[15:0]    reg_psum1_27_2;
wire[15:0]    reg_weight1_28_1;
wire[15:0]    reg_psum1_28_1;
wire[15:0]    reg_weight1_28_2;
wire[15:0]    reg_psum1_28_2;
wire[15:0]    reg_weight1_29_1;
wire[15:0]    reg_psum1_29_1;
wire[15:0]    reg_weight1_29_2;
wire[15:0]    reg_psum1_29_2;
wire[15:0]    reg_weight1_30_1;
wire[15:0]    reg_psum1_30_1;
wire[15:0]    reg_weight1_30_2;
wire[15:0]    reg_psum1_30_2;
wire[15:0]    reg_weight1_31_1;
wire[15:0]    reg_psum1_31_1;
wire[15:0]    reg_weight1_31_2;
wire[15:0]    reg_psum1_31_2;
wire[15:0]    reg_weight1_32_1;
wire[15:0]    reg_psum1_32_1;
wire[15:0]    reg_weight1_32_2;
wire[15:0]    reg_psum1_32_2;
wire[15:0]    reg_weight2_1_1;
wire[15:0]    reg_psum2_1_1;
wire[15:0]    reg_weight2_1_2;
wire[15:0]    reg_psum2_1_2;
wire[15:0]    reg_weight2_2_1;
wire[15:0]    reg_psum2_2_1;
wire[15:0]    reg_weight2_2_2;
wire[15:0]    reg_psum2_2_2;
wire[15:0]    reg_weight2_3_1;
wire[15:0]    reg_psum2_3_1;
wire[15:0]    reg_weight2_3_2;
wire[15:0]    reg_psum2_3_2;
wire[15:0]    reg_weight2_4_1;
wire[15:0]    reg_psum2_4_1;
wire[15:0]    reg_weight2_4_2;
wire[15:0]    reg_psum2_4_2;
wire[15:0]    reg_weight2_5_1;
wire[15:0]    reg_psum2_5_1;
wire[15:0]    reg_weight2_5_2;
wire[15:0]    reg_psum2_5_2;
wire[15:0]    reg_weight2_6_1;
wire[15:0]    reg_psum2_6_1;
wire[15:0]    reg_weight2_6_2;
wire[15:0]    reg_psum2_6_2;
wire[15:0]    reg_weight2_7_1;
wire[15:0]    reg_psum2_7_1;
wire[15:0]    reg_weight2_7_2;
wire[15:0]    reg_psum2_7_2;
wire[15:0]    reg_weight2_8_1;
wire[15:0]    reg_psum2_8_1;
wire[15:0]    reg_weight2_8_2;
wire[15:0]    reg_psum2_8_2;
wire[15:0]    reg_weight2_9_1;
wire[15:0]    reg_psum2_9_1;
wire[15:0]    reg_weight2_9_2;
wire[15:0]    reg_psum2_9_2;
wire[15:0]    reg_weight2_10_1;
wire[15:0]    reg_psum2_10_1;
wire[15:0]    reg_weight2_10_2;
wire[15:0]    reg_psum2_10_2;
wire[15:0]    reg_weight2_11_1;
wire[15:0]    reg_psum2_11_1;
wire[15:0]    reg_weight2_11_2;
wire[15:0]    reg_psum2_11_2;
wire[15:0]    reg_weight2_12_1;
wire[15:0]    reg_psum2_12_1;
wire[15:0]    reg_weight2_12_2;
wire[15:0]    reg_psum2_12_2;
wire[15:0]    reg_weight2_13_1;
wire[15:0]    reg_psum2_13_1;
wire[15:0]    reg_weight2_13_2;
wire[15:0]    reg_psum2_13_2;
wire[15:0]    reg_weight2_14_1;
wire[15:0]    reg_psum2_14_1;
wire[15:0]    reg_weight2_14_2;
wire[15:0]    reg_psum2_14_2;
wire[15:0]    reg_weight2_15_1;
wire[15:0]    reg_psum2_15_1;
wire[15:0]    reg_weight2_15_2;
wire[15:0]    reg_psum2_15_2;
wire[15:0]    reg_weight2_16_1;
wire[15:0]    reg_psum2_16_1;
wire[15:0]    reg_weight2_16_2;
wire[15:0]    reg_psum2_16_2;
wire[15:0]    reg_weight2_17_1;
wire[15:0]    reg_psum2_17_1;
wire[15:0]    reg_weight2_17_2;
wire[15:0]    reg_psum2_17_2;
wire[15:0]    reg_weight2_18_1;
wire[15:0]    reg_psum2_18_1;
wire[15:0]    reg_weight2_18_2;
wire[15:0]    reg_psum2_18_2;
wire[15:0]    reg_weight2_19_1;
wire[15:0]    reg_psum2_19_1;
wire[15:0]    reg_weight2_19_2;
wire[15:0]    reg_psum2_19_2;
wire[15:0]    reg_weight2_20_1;
wire[15:0]    reg_psum2_20_1;
wire[15:0]    reg_weight2_20_2;
wire[15:0]    reg_psum2_20_2;
wire[15:0]    reg_weight2_21_1;
wire[15:0]    reg_psum2_21_1;
wire[15:0]    reg_weight2_21_2;
wire[15:0]    reg_psum2_21_2;
wire[15:0]    reg_weight2_22_1;
wire[15:0]    reg_psum2_22_1;
wire[15:0]    reg_weight2_22_2;
wire[15:0]    reg_psum2_22_2;
wire[15:0]    reg_weight2_23_1;
wire[15:0]    reg_psum2_23_1;
wire[15:0]    reg_weight2_23_2;
wire[15:0]    reg_psum2_23_2;
wire[15:0]    reg_weight2_24_1;
wire[15:0]    reg_psum2_24_1;
wire[15:0]    reg_weight2_24_2;
wire[15:0]    reg_psum2_24_2;
wire[15:0]    reg_weight2_25_1;
wire[15:0]    reg_psum2_25_1;
wire[15:0]    reg_weight2_25_2;
wire[15:0]    reg_psum2_25_2;
wire[15:0]    reg_weight2_26_1;
wire[15:0]    reg_psum2_26_1;
wire[15:0]    reg_weight2_26_2;
wire[15:0]    reg_psum2_26_2;
wire[15:0]    reg_weight2_27_1;
wire[15:0]    reg_psum2_27_1;
wire[15:0]    reg_weight2_27_2;
wire[15:0]    reg_psum2_27_2;
wire[15:0]    reg_weight2_28_1;
wire[15:0]    reg_psum2_28_1;
wire[15:0]    reg_weight2_28_2;
wire[15:0]    reg_psum2_28_2;
wire[15:0]    reg_weight2_29_1;
wire[15:0]    reg_psum2_29_1;
wire[15:0]    reg_weight2_29_2;
wire[15:0]    reg_psum2_29_2;
wire[15:0]    reg_weight2_30_1;
wire[15:0]    reg_psum2_30_1;
wire[15:0]    reg_weight2_30_2;
wire[15:0]    reg_psum2_30_2;
wire[15:0]    reg_weight2_31_1;
wire[15:0]    reg_psum2_31_1;
wire[15:0]    reg_weight2_31_2;
wire[15:0]    reg_psum2_31_2;
wire[15:0]    reg_weight2_32_1;
wire[15:0]    reg_psum2_32_1;
wire[15:0]    reg_weight2_32_2;
wire[15:0]    reg_psum2_32_2;
wire[15:0]    reg_weight3_1_1;
wire[15:0]    reg_psum3_1_1;
wire[15:0]    reg_weight3_1_2;
wire[15:0]    reg_psum3_1_2;
wire[15:0]    reg_weight3_2_1;
wire[15:0]    reg_psum3_2_1;
wire[15:0]    reg_weight3_2_2;
wire[15:0]    reg_psum3_2_2;
wire[15:0]    reg_weight3_3_1;
wire[15:0]    reg_psum3_3_1;
wire[15:0]    reg_weight3_3_2;
wire[15:0]    reg_psum3_3_2;
wire[15:0]    reg_weight3_4_1;
wire[15:0]    reg_psum3_4_1;
wire[15:0]    reg_weight3_4_2;
wire[15:0]    reg_psum3_4_2;
wire[15:0]    reg_weight3_5_1;
wire[15:0]    reg_psum3_5_1;
wire[15:0]    reg_weight3_5_2;
wire[15:0]    reg_psum3_5_2;
wire[15:0]    reg_weight3_6_1;
wire[15:0]    reg_psum3_6_1;
wire[15:0]    reg_weight3_6_2;
wire[15:0]    reg_psum3_6_2;
wire[15:0]    reg_weight3_7_1;
wire[15:0]    reg_psum3_7_1;
wire[15:0]    reg_weight3_7_2;
wire[15:0]    reg_psum3_7_2;
wire[15:0]    reg_weight3_8_1;
wire[15:0]    reg_psum3_8_1;
wire[15:0]    reg_weight3_8_2;
wire[15:0]    reg_psum3_8_2;
wire[15:0]    reg_weight3_9_1;
wire[15:0]    reg_psum3_9_1;
wire[15:0]    reg_weight3_9_2;
wire[15:0]    reg_psum3_9_2;
wire[15:0]    reg_weight3_10_1;
wire[15:0]    reg_psum3_10_1;
wire[15:0]    reg_weight3_10_2;
wire[15:0]    reg_psum3_10_2;
wire[15:0]    reg_weight3_11_1;
wire[15:0]    reg_psum3_11_1;
wire[15:0]    reg_weight3_11_2;
wire[15:0]    reg_psum3_11_2;
wire[15:0]    reg_weight3_12_1;
wire[15:0]    reg_psum3_12_1;
wire[15:0]    reg_weight3_12_2;
wire[15:0]    reg_psum3_12_2;
wire[15:0]    reg_weight3_13_1;
wire[15:0]    reg_psum3_13_1;
wire[15:0]    reg_weight3_13_2;
wire[15:0]    reg_psum3_13_2;
wire[15:0]    reg_weight3_14_1;
wire[15:0]    reg_psum3_14_1;
wire[15:0]    reg_weight3_14_2;
wire[15:0]    reg_psum3_14_2;
wire[15:0]    reg_weight3_15_1;
wire[15:0]    reg_psum3_15_1;
wire[15:0]    reg_weight3_15_2;
wire[15:0]    reg_psum3_15_2;
wire[15:0]    reg_weight3_16_1;
wire[15:0]    reg_psum3_16_1;
wire[15:0]    reg_weight3_16_2;
wire[15:0]    reg_psum3_16_2;
wire[15:0]    reg_weight3_17_1;
wire[15:0]    reg_psum3_17_1;
wire[15:0]    reg_weight3_17_2;
wire[15:0]    reg_psum3_17_2;
wire[15:0]    reg_weight3_18_1;
wire[15:0]    reg_psum3_18_1;
wire[15:0]    reg_weight3_18_2;
wire[15:0]    reg_psum3_18_2;
wire[15:0]    reg_weight3_19_1;
wire[15:0]    reg_psum3_19_1;
wire[15:0]    reg_weight3_19_2;
wire[15:0]    reg_psum3_19_2;
wire[15:0]    reg_weight3_20_1;
wire[15:0]    reg_psum3_20_1;
wire[15:0]    reg_weight3_20_2;
wire[15:0]    reg_psum3_20_2;
wire[15:0]    reg_weight3_21_1;
wire[15:0]    reg_psum3_21_1;
wire[15:0]    reg_weight3_21_2;
wire[15:0]    reg_psum3_21_2;
wire[15:0]    reg_weight3_22_1;
wire[15:0]    reg_psum3_22_1;
wire[15:0]    reg_weight3_22_2;
wire[15:0]    reg_psum3_22_2;
wire[15:0]    reg_weight3_23_1;
wire[15:0]    reg_psum3_23_1;
wire[15:0]    reg_weight3_23_2;
wire[15:0]    reg_psum3_23_2;
wire[15:0]    reg_weight3_24_1;
wire[15:0]    reg_psum3_24_1;
wire[15:0]    reg_weight3_24_2;
wire[15:0]    reg_psum3_24_2;
wire[15:0]    reg_weight3_25_1;
wire[15:0]    reg_psum3_25_1;
wire[15:0]    reg_weight3_25_2;
wire[15:0]    reg_psum3_25_2;
wire[15:0]    reg_weight3_26_1;
wire[15:0]    reg_psum3_26_1;
wire[15:0]    reg_weight3_26_2;
wire[15:0]    reg_psum3_26_2;
wire[15:0]    reg_weight3_27_1;
wire[15:0]    reg_psum3_27_1;
wire[15:0]    reg_weight3_27_2;
wire[15:0]    reg_psum3_27_2;
wire[15:0]    reg_weight3_28_1;
wire[15:0]    reg_psum3_28_1;
wire[15:0]    reg_weight3_28_2;
wire[15:0]    reg_psum3_28_2;
wire[15:0]    reg_weight3_29_1;
wire[15:0]    reg_psum3_29_1;
wire[15:0]    reg_weight3_29_2;
wire[15:0]    reg_psum3_29_2;
wire[15:0]    reg_weight3_30_1;
wire[15:0]    reg_psum3_30_1;
wire[15:0]    reg_weight3_30_2;
wire[15:0]    reg_psum3_30_2;
wire[15:0]    reg_weight3_31_1;
wire[15:0]    reg_psum3_31_1;
wire[15:0]    reg_weight3_31_2;
wire[15:0]    reg_psum3_31_2;
wire[15:0]    reg_weight3_32_1;
wire[15:0]    reg_psum3_32_1;
wire[15:0]    reg_weight3_32_2;
wire[15:0]    reg_psum3_32_2;
wire[15:0]    reg_weight4_1_1;
wire[15:0]    reg_psum4_1_1;
wire[15:0]    reg_weight4_1_2;
wire[15:0]    reg_psum4_1_2;
wire[15:0]    reg_weight4_2_1;
wire[15:0]    reg_psum4_2_1;
wire[15:0]    reg_weight4_2_2;
wire[15:0]    reg_psum4_2_2;
wire[15:0]    reg_weight4_3_1;
wire[15:0]    reg_psum4_3_1;
wire[15:0]    reg_weight4_3_2;
wire[15:0]    reg_psum4_3_2;
wire[15:0]    reg_weight4_4_1;
wire[15:0]    reg_psum4_4_1;
wire[15:0]    reg_weight4_4_2;
wire[15:0]    reg_psum4_4_2;
wire[15:0]    reg_weight4_5_1;
wire[15:0]    reg_psum4_5_1;
wire[15:0]    reg_weight4_5_2;
wire[15:0]    reg_psum4_5_2;
wire[15:0]    reg_weight4_6_1;
wire[15:0]    reg_psum4_6_1;
wire[15:0]    reg_weight4_6_2;
wire[15:0]    reg_psum4_6_2;
wire[15:0]    reg_weight4_7_1;
wire[15:0]    reg_psum4_7_1;
wire[15:0]    reg_weight4_7_2;
wire[15:0]    reg_psum4_7_2;
wire[15:0]    reg_weight4_8_1;
wire[15:0]    reg_psum4_8_1;
wire[15:0]    reg_weight4_8_2;
wire[15:0]    reg_psum4_8_2;
wire[15:0]    reg_weight4_9_1;
wire[15:0]    reg_psum4_9_1;
wire[15:0]    reg_weight4_9_2;
wire[15:0]    reg_psum4_9_2;
wire[15:0]    reg_weight4_10_1;
wire[15:0]    reg_psum4_10_1;
wire[15:0]    reg_weight4_10_2;
wire[15:0]    reg_psum4_10_2;
wire[15:0]    reg_weight4_11_1;
wire[15:0]    reg_psum4_11_1;
wire[15:0]    reg_weight4_11_2;
wire[15:0]    reg_psum4_11_2;
wire[15:0]    reg_weight4_12_1;
wire[15:0]    reg_psum4_12_1;
wire[15:0]    reg_weight4_12_2;
wire[15:0]    reg_psum4_12_2;
wire[15:0]    reg_weight4_13_1;
wire[15:0]    reg_psum4_13_1;
wire[15:0]    reg_weight4_13_2;
wire[15:0]    reg_psum4_13_2;
wire[15:0]    reg_weight4_14_1;
wire[15:0]    reg_psum4_14_1;
wire[15:0]    reg_weight4_14_2;
wire[15:0]    reg_psum4_14_2;
wire[15:0]    reg_weight4_15_1;
wire[15:0]    reg_psum4_15_1;
wire[15:0]    reg_weight4_15_2;
wire[15:0]    reg_psum4_15_2;
wire[15:0]    reg_weight4_16_1;
wire[15:0]    reg_psum4_16_1;
wire[15:0]    reg_weight4_16_2;
wire[15:0]    reg_psum4_16_2;
wire[15:0]    reg_weight4_17_1;
wire[15:0]    reg_psum4_17_1;
wire[15:0]    reg_weight4_17_2;
wire[15:0]    reg_psum4_17_2;
wire[15:0]    reg_weight4_18_1;
wire[15:0]    reg_psum4_18_1;
wire[15:0]    reg_weight4_18_2;
wire[15:0]    reg_psum4_18_2;
wire[15:0]    reg_weight4_19_1;
wire[15:0]    reg_psum4_19_1;
wire[15:0]    reg_weight4_19_2;
wire[15:0]    reg_psum4_19_2;
wire[15:0]    reg_weight4_20_1;
wire[15:0]    reg_psum4_20_1;
wire[15:0]    reg_weight4_20_2;
wire[15:0]    reg_psum4_20_2;
wire[15:0]    reg_weight4_21_1;
wire[15:0]    reg_psum4_21_1;
wire[15:0]    reg_weight4_21_2;
wire[15:0]    reg_psum4_21_2;
wire[15:0]    reg_weight4_22_1;
wire[15:0]    reg_psum4_22_1;
wire[15:0]    reg_weight4_22_2;
wire[15:0]    reg_psum4_22_2;
wire[15:0]    reg_weight4_23_1;
wire[15:0]    reg_psum4_23_1;
wire[15:0]    reg_weight4_23_2;
wire[15:0]    reg_psum4_23_2;
wire[15:0]    reg_weight4_24_1;
wire[15:0]    reg_psum4_24_1;
wire[15:0]    reg_weight4_24_2;
wire[15:0]    reg_psum4_24_2;
wire[15:0]    reg_weight4_25_1;
wire[15:0]    reg_psum4_25_1;
wire[15:0]    reg_weight4_25_2;
wire[15:0]    reg_psum4_25_2;
wire[15:0]    reg_weight4_26_1;
wire[15:0]    reg_psum4_26_1;
wire[15:0]    reg_weight4_26_2;
wire[15:0]    reg_psum4_26_2;
wire[15:0]    reg_weight4_27_1;
wire[15:0]    reg_psum4_27_1;
wire[15:0]    reg_weight4_27_2;
wire[15:0]    reg_psum4_27_2;
wire[15:0]    reg_weight4_28_1;
wire[15:0]    reg_psum4_28_1;
wire[15:0]    reg_weight4_28_2;
wire[15:0]    reg_psum4_28_2;
wire[15:0]    reg_weight4_29_1;
wire[15:0]    reg_psum4_29_1;
wire[15:0]    reg_weight4_29_2;
wire[15:0]    reg_psum4_29_2;
wire[15:0]    reg_weight4_30_1;
wire[15:0]    reg_psum4_30_1;
wire[15:0]    reg_weight4_30_2;
wire[15:0]    reg_psum4_30_2;
wire[15:0]    reg_weight4_31_1;
wire[15:0]    reg_psum4_31_1;
wire[15:0]    reg_weight4_31_2;
wire[15:0]    reg_psum4_31_2;
wire[15:0]    reg_weight4_32_1;
wire[15:0]    reg_psum4_32_1;
wire[15:0]    reg_weight4_32_2;
wire[15:0]    reg_psum4_32_2;
wire[15:0]    reg_weight5_1_1;
wire[15:0]    reg_psum5_1_1;
wire[15:0]    reg_weight5_1_2;
wire[15:0]    reg_psum5_1_2;
wire[15:0]    reg_weight5_2_1;
wire[15:0]    reg_psum5_2_1;
wire[15:0]    reg_weight5_2_2;
wire[15:0]    reg_psum5_2_2;
wire[15:0]    reg_weight5_3_1;
wire[15:0]    reg_psum5_3_1;
wire[15:0]    reg_weight5_3_2;
wire[15:0]    reg_psum5_3_2;
wire[15:0]    reg_weight5_4_1;
wire[15:0]    reg_psum5_4_1;
wire[15:0]    reg_weight5_4_2;
wire[15:0]    reg_psum5_4_2;
wire[15:0]    reg_weight5_5_1;
wire[15:0]    reg_psum5_5_1;
wire[15:0]    reg_weight5_5_2;
wire[15:0]    reg_psum5_5_2;
wire[15:0]    reg_weight5_6_1;
wire[15:0]    reg_psum5_6_1;
wire[15:0]    reg_weight5_6_2;
wire[15:0]    reg_psum5_6_2;
wire[15:0]    reg_weight5_7_1;
wire[15:0]    reg_psum5_7_1;
wire[15:0]    reg_weight5_7_2;
wire[15:0]    reg_psum5_7_2;
wire[15:0]    reg_weight5_8_1;
wire[15:0]    reg_psum5_8_1;
wire[15:0]    reg_weight5_8_2;
wire[15:0]    reg_psum5_8_2;
wire[15:0]    reg_weight5_9_1;
wire[15:0]    reg_psum5_9_1;
wire[15:0]    reg_weight5_9_2;
wire[15:0]    reg_psum5_9_2;
wire[15:0]    reg_weight5_10_1;
wire[15:0]    reg_psum5_10_1;
wire[15:0]    reg_weight5_10_2;
wire[15:0]    reg_psum5_10_2;
wire[15:0]    reg_weight5_11_1;
wire[15:0]    reg_psum5_11_1;
wire[15:0]    reg_weight5_11_2;
wire[15:0]    reg_psum5_11_2;
wire[15:0]    reg_weight5_12_1;
wire[15:0]    reg_psum5_12_1;
wire[15:0]    reg_weight5_12_2;
wire[15:0]    reg_psum5_12_2;
wire[15:0]    reg_weight5_13_1;
wire[15:0]    reg_psum5_13_1;
wire[15:0]    reg_weight5_13_2;
wire[15:0]    reg_psum5_13_2;
wire[15:0]    reg_weight5_14_1;
wire[15:0]    reg_psum5_14_1;
wire[15:0]    reg_weight5_14_2;
wire[15:0]    reg_psum5_14_2;
wire[15:0]    reg_weight5_15_1;
wire[15:0]    reg_psum5_15_1;
wire[15:0]    reg_weight5_15_2;
wire[15:0]    reg_psum5_15_2;
wire[15:0]    reg_weight5_16_1;
wire[15:0]    reg_psum5_16_1;
wire[15:0]    reg_weight5_16_2;
wire[15:0]    reg_psum5_16_2;
wire[15:0]    reg_weight5_17_1;
wire[15:0]    reg_psum5_17_1;
wire[15:0]    reg_weight5_17_2;
wire[15:0]    reg_psum5_17_2;
wire[15:0]    reg_weight5_18_1;
wire[15:0]    reg_psum5_18_1;
wire[15:0]    reg_weight5_18_2;
wire[15:0]    reg_psum5_18_2;
wire[15:0]    reg_weight5_19_1;
wire[15:0]    reg_psum5_19_1;
wire[15:0]    reg_weight5_19_2;
wire[15:0]    reg_psum5_19_2;
wire[15:0]    reg_weight5_20_1;
wire[15:0]    reg_psum5_20_1;
wire[15:0]    reg_weight5_20_2;
wire[15:0]    reg_psum5_20_2;
wire[15:0]    reg_weight5_21_1;
wire[15:0]    reg_psum5_21_1;
wire[15:0]    reg_weight5_21_2;
wire[15:0]    reg_psum5_21_2;
wire[15:0]    reg_weight5_22_1;
wire[15:0]    reg_psum5_22_1;
wire[15:0]    reg_weight5_22_2;
wire[15:0]    reg_psum5_22_2;
wire[15:0]    reg_weight5_23_1;
wire[15:0]    reg_psum5_23_1;
wire[15:0]    reg_weight5_23_2;
wire[15:0]    reg_psum5_23_2;
wire[15:0]    reg_weight5_24_1;
wire[15:0]    reg_psum5_24_1;
wire[15:0]    reg_weight5_24_2;
wire[15:0]    reg_psum5_24_2;
wire[15:0]    reg_weight5_25_1;
wire[15:0]    reg_psum5_25_1;
wire[15:0]    reg_weight5_25_2;
wire[15:0]    reg_psum5_25_2;
wire[15:0]    reg_weight5_26_1;
wire[15:0]    reg_psum5_26_1;
wire[15:0]    reg_weight5_26_2;
wire[15:0]    reg_psum5_26_2;
wire[15:0]    reg_weight5_27_1;
wire[15:0]    reg_psum5_27_1;
wire[15:0]    reg_weight5_27_2;
wire[15:0]    reg_psum5_27_2;
wire[15:0]    reg_weight5_28_1;
wire[15:0]    reg_psum5_28_1;
wire[15:0]    reg_weight5_28_2;
wire[15:0]    reg_psum5_28_2;
wire[15:0]    reg_weight5_29_1;
wire[15:0]    reg_psum5_29_1;
wire[15:0]    reg_weight5_29_2;
wire[15:0]    reg_psum5_29_2;
wire[15:0]    reg_weight5_30_1;
wire[15:0]    reg_psum5_30_1;
wire[15:0]    reg_weight5_30_2;
wire[15:0]    reg_psum5_30_2;
wire[15:0]    reg_weight5_31_1;
wire[15:0]    reg_psum5_31_1;
wire[15:0]    reg_weight5_31_2;
wire[15:0]    reg_psum5_31_2;
wire[15:0]    reg_weight5_32_1;
wire[15:0]    reg_psum5_32_1;
wire[15:0]    reg_weight5_32_2;
wire[15:0]    reg_psum5_32_2;
wire[15:0]    reg_weight6_1_1;
wire[15:0]    reg_psum6_1_1;
wire[15:0]    reg_weight6_1_2;
wire[15:0]    reg_psum6_1_2;
wire[15:0]    reg_weight6_2_1;
wire[15:0]    reg_psum6_2_1;
wire[15:0]    reg_weight6_2_2;
wire[15:0]    reg_psum6_2_2;
wire[15:0]    reg_weight6_3_1;
wire[15:0]    reg_psum6_3_1;
wire[15:0]    reg_weight6_3_2;
wire[15:0]    reg_psum6_3_2;
wire[15:0]    reg_weight6_4_1;
wire[15:0]    reg_psum6_4_1;
wire[15:0]    reg_weight6_4_2;
wire[15:0]    reg_psum6_4_2;
wire[15:0]    reg_weight6_5_1;
wire[15:0]    reg_psum6_5_1;
wire[15:0]    reg_weight6_5_2;
wire[15:0]    reg_psum6_5_2;
wire[15:0]    reg_weight6_6_1;
wire[15:0]    reg_psum6_6_1;
wire[15:0]    reg_weight6_6_2;
wire[15:0]    reg_psum6_6_2;
wire[15:0]    reg_weight6_7_1;
wire[15:0]    reg_psum6_7_1;
wire[15:0]    reg_weight6_7_2;
wire[15:0]    reg_psum6_7_2;
wire[15:0]    reg_weight6_8_1;
wire[15:0]    reg_psum6_8_1;
wire[15:0]    reg_weight6_8_2;
wire[15:0]    reg_psum6_8_2;
wire[15:0]    reg_weight6_9_1;
wire[15:0]    reg_psum6_9_1;
wire[15:0]    reg_weight6_9_2;
wire[15:0]    reg_psum6_9_2;
wire[15:0]    reg_weight6_10_1;
wire[15:0]    reg_psum6_10_1;
wire[15:0]    reg_weight6_10_2;
wire[15:0]    reg_psum6_10_2;
wire[15:0]    reg_weight6_11_1;
wire[15:0]    reg_psum6_11_1;
wire[15:0]    reg_weight6_11_2;
wire[15:0]    reg_psum6_11_2;
wire[15:0]    reg_weight6_12_1;
wire[15:0]    reg_psum6_12_1;
wire[15:0]    reg_weight6_12_2;
wire[15:0]    reg_psum6_12_2;
wire[15:0]    reg_weight6_13_1;
wire[15:0]    reg_psum6_13_1;
wire[15:0]    reg_weight6_13_2;
wire[15:0]    reg_psum6_13_2;
wire[15:0]    reg_weight6_14_1;
wire[15:0]    reg_psum6_14_1;
wire[15:0]    reg_weight6_14_2;
wire[15:0]    reg_psum6_14_2;
wire[15:0]    reg_weight6_15_1;
wire[15:0]    reg_psum6_15_1;
wire[15:0]    reg_weight6_15_2;
wire[15:0]    reg_psum6_15_2;
wire[15:0]    reg_weight6_16_1;
wire[15:0]    reg_psum6_16_1;
wire[15:0]    reg_weight6_16_2;
wire[15:0]    reg_psum6_16_2;
wire[15:0]    reg_weight6_17_1;
wire[15:0]    reg_psum6_17_1;
wire[15:0]    reg_weight6_17_2;
wire[15:0]    reg_psum6_17_2;
wire[15:0]    reg_weight6_18_1;
wire[15:0]    reg_psum6_18_1;
wire[15:0]    reg_weight6_18_2;
wire[15:0]    reg_psum6_18_2;
wire[15:0]    reg_weight6_19_1;
wire[15:0]    reg_psum6_19_1;
wire[15:0]    reg_weight6_19_2;
wire[15:0]    reg_psum6_19_2;
wire[15:0]    reg_weight6_20_1;
wire[15:0]    reg_psum6_20_1;
wire[15:0]    reg_weight6_20_2;
wire[15:0]    reg_psum6_20_2;
wire[15:0]    reg_weight6_21_1;
wire[15:0]    reg_psum6_21_1;
wire[15:0]    reg_weight6_21_2;
wire[15:0]    reg_psum6_21_2;
wire[15:0]    reg_weight6_22_1;
wire[15:0]    reg_psum6_22_1;
wire[15:0]    reg_weight6_22_2;
wire[15:0]    reg_psum6_22_2;
wire[15:0]    reg_weight6_23_1;
wire[15:0]    reg_psum6_23_1;
wire[15:0]    reg_weight6_23_2;
wire[15:0]    reg_psum6_23_2;
wire[15:0]    reg_weight6_24_1;
wire[15:0]    reg_psum6_24_1;
wire[15:0]    reg_weight6_24_2;
wire[15:0]    reg_psum6_24_2;
wire[15:0]    reg_weight6_25_1;
wire[15:0]    reg_psum6_25_1;
wire[15:0]    reg_weight6_25_2;
wire[15:0]    reg_psum6_25_2;
wire[15:0]    reg_weight6_26_1;
wire[15:0]    reg_psum6_26_1;
wire[15:0]    reg_weight6_26_2;
wire[15:0]    reg_psum6_26_2;
wire[15:0]    reg_weight6_27_1;
wire[15:0]    reg_psum6_27_1;
wire[15:0]    reg_weight6_27_2;
wire[15:0]    reg_psum6_27_2;
wire[15:0]    reg_weight6_28_1;
wire[15:0]    reg_psum6_28_1;
wire[15:0]    reg_weight6_28_2;
wire[15:0]    reg_psum6_28_2;
wire[15:0]    reg_weight6_29_1;
wire[15:0]    reg_psum6_29_1;
wire[15:0]    reg_weight6_29_2;
wire[15:0]    reg_psum6_29_2;
wire[15:0]    reg_weight6_30_1;
wire[15:0]    reg_psum6_30_1;
wire[15:0]    reg_weight6_30_2;
wire[15:0]    reg_psum6_30_2;
wire[15:0]    reg_weight6_31_1;
wire[15:0]    reg_psum6_31_1;
wire[15:0]    reg_weight6_31_2;
wire[15:0]    reg_psum6_31_2;
wire[15:0]    reg_weight6_32_1;
wire[15:0]    reg_psum6_32_1;
wire[15:0]    reg_weight6_32_2;
wire[15:0]    reg_psum6_32_2;
wire[15:0]    reg_weight7_1_1;
wire[15:0]    reg_psum7_1_1;
wire[15:0]    reg_weight7_1_2;
wire[15:0]    reg_psum7_1_2;
wire[15:0]    reg_weight7_2_1;
wire[15:0]    reg_psum7_2_1;
wire[15:0]    reg_weight7_2_2;
wire[15:0]    reg_psum7_2_2;
wire[15:0]    reg_weight7_3_1;
wire[15:0]    reg_psum7_3_1;
wire[15:0]    reg_weight7_3_2;
wire[15:0]    reg_psum7_3_2;
wire[15:0]    reg_weight7_4_1;
wire[15:0]    reg_psum7_4_1;
wire[15:0]    reg_weight7_4_2;
wire[15:0]    reg_psum7_4_2;
wire[15:0]    reg_weight7_5_1;
wire[15:0]    reg_psum7_5_1;
wire[15:0]    reg_weight7_5_2;
wire[15:0]    reg_psum7_5_2;
wire[15:0]    reg_weight7_6_1;
wire[15:0]    reg_psum7_6_1;
wire[15:0]    reg_weight7_6_2;
wire[15:0]    reg_psum7_6_2;
wire[15:0]    reg_weight7_7_1;
wire[15:0]    reg_psum7_7_1;
wire[15:0]    reg_weight7_7_2;
wire[15:0]    reg_psum7_7_2;
wire[15:0]    reg_weight7_8_1;
wire[15:0]    reg_psum7_8_1;
wire[15:0]    reg_weight7_8_2;
wire[15:0]    reg_psum7_8_2;
wire[15:0]    reg_weight7_9_1;
wire[15:0]    reg_psum7_9_1;
wire[15:0]    reg_weight7_9_2;
wire[15:0]    reg_psum7_9_2;
wire[15:0]    reg_weight7_10_1;
wire[15:0]    reg_psum7_10_1;
wire[15:0]    reg_weight7_10_2;
wire[15:0]    reg_psum7_10_2;
wire[15:0]    reg_weight7_11_1;
wire[15:0]    reg_psum7_11_1;
wire[15:0]    reg_weight7_11_2;
wire[15:0]    reg_psum7_11_2;
wire[15:0]    reg_weight7_12_1;
wire[15:0]    reg_psum7_12_1;
wire[15:0]    reg_weight7_12_2;
wire[15:0]    reg_psum7_12_2;
wire[15:0]    reg_weight7_13_1;
wire[15:0]    reg_psum7_13_1;
wire[15:0]    reg_weight7_13_2;
wire[15:0]    reg_psum7_13_2;
wire[15:0]    reg_weight7_14_1;
wire[15:0]    reg_psum7_14_1;
wire[15:0]    reg_weight7_14_2;
wire[15:0]    reg_psum7_14_2;
wire[15:0]    reg_weight7_15_1;
wire[15:0]    reg_psum7_15_1;
wire[15:0]    reg_weight7_15_2;
wire[15:0]    reg_psum7_15_2;
wire[15:0]    reg_weight7_16_1;
wire[15:0]    reg_psum7_16_1;
wire[15:0]    reg_weight7_16_2;
wire[15:0]    reg_psum7_16_2;
wire[15:0]    reg_weight7_17_1;
wire[15:0]    reg_psum7_17_1;
wire[15:0]    reg_weight7_17_2;
wire[15:0]    reg_psum7_17_2;
wire[15:0]    reg_weight7_18_1;
wire[15:0]    reg_psum7_18_1;
wire[15:0]    reg_weight7_18_2;
wire[15:0]    reg_psum7_18_2;
wire[15:0]    reg_weight7_19_1;
wire[15:0]    reg_psum7_19_1;
wire[15:0]    reg_weight7_19_2;
wire[15:0]    reg_psum7_19_2;
wire[15:0]    reg_weight7_20_1;
wire[15:0]    reg_psum7_20_1;
wire[15:0]    reg_weight7_20_2;
wire[15:0]    reg_psum7_20_2;
wire[15:0]    reg_weight7_21_1;
wire[15:0]    reg_psum7_21_1;
wire[15:0]    reg_weight7_21_2;
wire[15:0]    reg_psum7_21_2;
wire[15:0]    reg_weight7_22_1;
wire[15:0]    reg_psum7_22_1;
wire[15:0]    reg_weight7_22_2;
wire[15:0]    reg_psum7_22_2;
wire[15:0]    reg_weight7_23_1;
wire[15:0]    reg_psum7_23_1;
wire[15:0]    reg_weight7_23_2;
wire[15:0]    reg_psum7_23_2;
wire[15:0]    reg_weight7_24_1;
wire[15:0]    reg_psum7_24_1;
wire[15:0]    reg_weight7_24_2;
wire[15:0]    reg_psum7_24_2;
wire[15:0]    reg_weight7_25_1;
wire[15:0]    reg_psum7_25_1;
wire[15:0]    reg_weight7_25_2;
wire[15:0]    reg_psum7_25_2;
wire[15:0]    reg_weight7_26_1;
wire[15:0]    reg_psum7_26_1;
wire[15:0]    reg_weight7_26_2;
wire[15:0]    reg_psum7_26_2;
wire[15:0]    reg_weight7_27_1;
wire[15:0]    reg_psum7_27_1;
wire[15:0]    reg_weight7_27_2;
wire[15:0]    reg_psum7_27_2;
wire[15:0]    reg_weight7_28_1;
wire[15:0]    reg_psum7_28_1;
wire[15:0]    reg_weight7_28_2;
wire[15:0]    reg_psum7_28_2;
wire[15:0]    reg_weight7_29_1;
wire[15:0]    reg_psum7_29_1;
wire[15:0]    reg_weight7_29_2;
wire[15:0]    reg_psum7_29_2;
wire[15:0]    reg_weight7_30_1;
wire[15:0]    reg_psum7_30_1;
wire[15:0]    reg_weight7_30_2;
wire[15:0]    reg_psum7_30_2;
wire[15:0]    reg_weight7_31_1;
wire[15:0]    reg_psum7_31_1;
wire[15:0]    reg_weight7_31_2;
wire[15:0]    reg_psum7_31_2;
wire[15:0]    reg_weight7_32_1;
wire[15:0]    reg_psum7_32_1;
wire[15:0]    reg_weight7_32_2;
wire[15:0]    reg_psum7_32_2;
wire[15:0]    reg_weight8_1_1;
wire[15:0]    reg_psum8_1_1;
wire[15:0]    reg_weight8_1_2;
wire[15:0]    reg_psum8_1_2;
wire[15:0]    reg_weight8_2_1;
wire[15:0]    reg_psum8_2_1;
wire[15:0]    reg_weight8_2_2;
wire[15:0]    reg_psum8_2_2;
wire[15:0]    reg_weight8_3_1;
wire[15:0]    reg_psum8_3_1;
wire[15:0]    reg_weight8_3_2;
wire[15:0]    reg_psum8_3_2;
wire[15:0]    reg_weight8_4_1;
wire[15:0]    reg_psum8_4_1;
wire[15:0]    reg_weight8_4_2;
wire[15:0]    reg_psum8_4_2;
wire[15:0]    reg_weight8_5_1;
wire[15:0]    reg_psum8_5_1;
wire[15:0]    reg_weight8_5_2;
wire[15:0]    reg_psum8_5_2;
wire[15:0]    reg_weight8_6_1;
wire[15:0]    reg_psum8_6_1;
wire[15:0]    reg_weight8_6_2;
wire[15:0]    reg_psum8_6_2;
wire[15:0]    reg_weight8_7_1;
wire[15:0]    reg_psum8_7_1;
wire[15:0]    reg_weight8_7_2;
wire[15:0]    reg_psum8_7_2;
wire[15:0]    reg_weight8_8_1;
wire[15:0]    reg_psum8_8_1;
wire[15:0]    reg_weight8_8_2;
wire[15:0]    reg_psum8_8_2;
wire[15:0]    reg_weight8_9_1;
wire[15:0]    reg_psum8_9_1;
wire[15:0]    reg_weight8_9_2;
wire[15:0]    reg_psum8_9_2;
wire[15:0]    reg_weight8_10_1;
wire[15:0]    reg_psum8_10_1;
wire[15:0]    reg_weight8_10_2;
wire[15:0]    reg_psum8_10_2;
wire[15:0]    reg_weight8_11_1;
wire[15:0]    reg_psum8_11_1;
wire[15:0]    reg_weight8_11_2;
wire[15:0]    reg_psum8_11_2;
wire[15:0]    reg_weight8_12_1;
wire[15:0]    reg_psum8_12_1;
wire[15:0]    reg_weight8_12_2;
wire[15:0]    reg_psum8_12_2;
wire[15:0]    reg_weight8_13_1;
wire[15:0]    reg_psum8_13_1;
wire[15:0]    reg_weight8_13_2;
wire[15:0]    reg_psum8_13_2;
wire[15:0]    reg_weight8_14_1;
wire[15:0]    reg_psum8_14_1;
wire[15:0]    reg_weight8_14_2;
wire[15:0]    reg_psum8_14_2;
wire[15:0]    reg_weight8_15_1;
wire[15:0]    reg_psum8_15_1;
wire[15:0]    reg_weight8_15_2;
wire[15:0]    reg_psum8_15_2;
wire[15:0]    reg_weight8_16_1;
wire[15:0]    reg_psum8_16_1;
wire[15:0]    reg_weight8_16_2;
wire[15:0]    reg_psum8_16_2;
wire[15:0]    reg_weight8_17_1;
wire[15:0]    reg_psum8_17_1;
wire[15:0]    reg_weight8_17_2;
wire[15:0]    reg_psum8_17_2;
wire[15:0]    reg_weight8_18_1;
wire[15:0]    reg_psum8_18_1;
wire[15:0]    reg_weight8_18_2;
wire[15:0]    reg_psum8_18_2;
wire[15:0]    reg_weight8_19_1;
wire[15:0]    reg_psum8_19_1;
wire[15:0]    reg_weight8_19_2;
wire[15:0]    reg_psum8_19_2;
wire[15:0]    reg_weight8_20_1;
wire[15:0]    reg_psum8_20_1;
wire[15:0]    reg_weight8_20_2;
wire[15:0]    reg_psum8_20_2;
wire[15:0]    reg_weight8_21_1;
wire[15:0]    reg_psum8_21_1;
wire[15:0]    reg_weight8_21_2;
wire[15:0]    reg_psum8_21_2;
wire[15:0]    reg_weight8_22_1;
wire[15:0]    reg_psum8_22_1;
wire[15:0]    reg_weight8_22_2;
wire[15:0]    reg_psum8_22_2;
wire[15:0]    reg_weight8_23_1;
wire[15:0]    reg_psum8_23_1;
wire[15:0]    reg_weight8_23_2;
wire[15:0]    reg_psum8_23_2;
wire[15:0]    reg_weight8_24_1;
wire[15:0]    reg_psum8_24_1;
wire[15:0]    reg_weight8_24_2;
wire[15:0]    reg_psum8_24_2;
wire[15:0]    reg_weight8_25_1;
wire[15:0]    reg_psum8_25_1;
wire[15:0]    reg_weight8_25_2;
wire[15:0]    reg_psum8_25_2;
wire[15:0]    reg_weight8_26_1;
wire[15:0]    reg_psum8_26_1;
wire[15:0]    reg_weight8_26_2;
wire[15:0]    reg_psum8_26_2;
wire[15:0]    reg_weight8_27_1;
wire[15:0]    reg_psum8_27_1;
wire[15:0]    reg_weight8_27_2;
wire[15:0]    reg_psum8_27_2;
wire[15:0]    reg_weight8_28_1;
wire[15:0]    reg_psum8_28_1;
wire[15:0]    reg_weight8_28_2;
wire[15:0]    reg_psum8_28_2;
wire[15:0]    reg_weight8_29_1;
wire[15:0]    reg_psum8_29_1;
wire[15:0]    reg_weight8_29_2;
wire[15:0]    reg_psum8_29_2;
wire[15:0]    reg_weight8_30_1;
wire[15:0]    reg_psum8_30_1;
wire[15:0]    reg_weight8_30_2;
wire[15:0]    reg_psum8_30_2;
wire[15:0]    reg_weight8_31_1;
wire[15:0]    reg_psum8_31_1;
wire[15:0]    reg_weight8_31_2;
wire[15:0]    reg_psum8_31_2;
wire[15:0]    reg_weight8_32_1;
wire[15:0]    reg_psum8_32_1;
wire[15:0]    reg_weight8_32_2;
wire[15:0]    reg_psum8_32_2;
wire[15:0]    reg_weight9_1_1;
wire[15:0]    reg_psum9_1_1;
wire[15:0]    reg_weight9_1_2;
wire[15:0]    reg_psum9_1_2;
wire[15:0]    reg_weight9_2_1;
wire[15:0]    reg_psum9_2_1;
wire[15:0]    reg_weight9_2_2;
wire[15:0]    reg_psum9_2_2;
wire[15:0]    reg_weight9_3_1;
wire[15:0]    reg_psum9_3_1;
wire[15:0]    reg_weight9_3_2;
wire[15:0]    reg_psum9_3_2;
wire[15:0]    reg_weight9_4_1;
wire[15:0]    reg_psum9_4_1;
wire[15:0]    reg_weight9_4_2;
wire[15:0]    reg_psum9_4_2;
wire[15:0]    reg_weight9_5_1;
wire[15:0]    reg_psum9_5_1;
wire[15:0]    reg_weight9_5_2;
wire[15:0]    reg_psum9_5_2;
wire[15:0]    reg_weight9_6_1;
wire[15:0]    reg_psum9_6_1;
wire[15:0]    reg_weight9_6_2;
wire[15:0]    reg_psum9_6_2;
wire[15:0]    reg_weight9_7_1;
wire[15:0]    reg_psum9_7_1;
wire[15:0]    reg_weight9_7_2;
wire[15:0]    reg_psum9_7_2;
wire[15:0]    reg_weight9_8_1;
wire[15:0]    reg_psum9_8_1;
wire[15:0]    reg_weight9_8_2;
wire[15:0]    reg_psum9_8_2;
wire[15:0]    reg_weight9_9_1;
wire[15:0]    reg_psum9_9_1;
wire[15:0]    reg_weight9_9_2;
wire[15:0]    reg_psum9_9_2;
wire[15:0]    reg_weight9_10_1;
wire[15:0]    reg_psum9_10_1;
wire[15:0]    reg_weight9_10_2;
wire[15:0]    reg_psum9_10_2;
wire[15:0]    reg_weight9_11_1;
wire[15:0]    reg_psum9_11_1;
wire[15:0]    reg_weight9_11_2;
wire[15:0]    reg_psum9_11_2;
wire[15:0]    reg_weight9_12_1;
wire[15:0]    reg_psum9_12_1;
wire[15:0]    reg_weight9_12_2;
wire[15:0]    reg_psum9_12_2;
wire[15:0]    reg_weight9_13_1;
wire[15:0]    reg_psum9_13_1;
wire[15:0]    reg_weight9_13_2;
wire[15:0]    reg_psum9_13_2;
wire[15:0]    reg_weight9_14_1;
wire[15:0]    reg_psum9_14_1;
wire[15:0]    reg_weight9_14_2;
wire[15:0]    reg_psum9_14_2;
wire[15:0]    reg_weight9_15_1;
wire[15:0]    reg_psum9_15_1;
wire[15:0]    reg_weight9_15_2;
wire[15:0]    reg_psum9_15_2;
wire[15:0]    reg_weight9_16_1;
wire[15:0]    reg_psum9_16_1;
wire[15:0]    reg_weight9_16_2;
wire[15:0]    reg_psum9_16_2;
wire[15:0]    reg_weight9_17_1;
wire[15:0]    reg_psum9_17_1;
wire[15:0]    reg_weight9_17_2;
wire[15:0]    reg_psum9_17_2;
wire[15:0]    reg_weight9_18_1;
wire[15:0]    reg_psum9_18_1;
wire[15:0]    reg_weight9_18_2;
wire[15:0]    reg_psum9_18_2;
wire[15:0]    reg_weight9_19_1;
wire[15:0]    reg_psum9_19_1;
wire[15:0]    reg_weight9_19_2;
wire[15:0]    reg_psum9_19_2;
wire[15:0]    reg_weight9_20_1;
wire[15:0]    reg_psum9_20_1;
wire[15:0]    reg_weight9_20_2;
wire[15:0]    reg_psum9_20_2;
wire[15:0]    reg_weight9_21_1;
wire[15:0]    reg_psum9_21_1;
wire[15:0]    reg_weight9_21_2;
wire[15:0]    reg_psum9_21_2;
wire[15:0]    reg_weight9_22_1;
wire[15:0]    reg_psum9_22_1;
wire[15:0]    reg_weight9_22_2;
wire[15:0]    reg_psum9_22_2;
wire[15:0]    reg_weight9_23_1;
wire[15:0]    reg_psum9_23_1;
wire[15:0]    reg_weight9_23_2;
wire[15:0]    reg_psum9_23_2;
wire[15:0]    reg_weight9_24_1;
wire[15:0]    reg_psum9_24_1;
wire[15:0]    reg_weight9_24_2;
wire[15:0]    reg_psum9_24_2;
wire[15:0]    reg_weight9_25_1;
wire[15:0]    reg_psum9_25_1;
wire[15:0]    reg_weight9_25_2;
wire[15:0]    reg_psum9_25_2;
wire[15:0]    reg_weight9_26_1;
wire[15:0]    reg_psum9_26_1;
wire[15:0]    reg_weight9_26_2;
wire[15:0]    reg_psum9_26_2;
wire[15:0]    reg_weight9_27_1;
wire[15:0]    reg_psum9_27_1;
wire[15:0]    reg_weight9_27_2;
wire[15:0]    reg_psum9_27_2;
wire[15:0]    reg_weight9_28_1;
wire[15:0]    reg_psum9_28_1;
wire[15:0]    reg_weight9_28_2;
wire[15:0]    reg_psum9_28_2;
wire[15:0]    reg_weight9_29_1;
wire[15:0]    reg_psum9_29_1;
wire[15:0]    reg_weight9_29_2;
wire[15:0]    reg_psum9_29_2;
wire[15:0]    reg_weight9_30_1;
wire[15:0]    reg_psum9_30_1;
wire[15:0]    reg_weight9_30_2;
wire[15:0]    reg_psum9_30_2;
wire[15:0]    reg_weight9_31_1;
wire[15:0]    reg_psum9_31_1;
wire[15:0]    reg_weight9_31_2;
wire[15:0]    reg_psum9_31_2;
wire[15:0]    reg_weight9_32_1;
wire[15:0]    reg_psum9_32_1;
wire[15:0]    reg_weight9_32_2;
wire[15:0]    reg_psum9_32_2;
wire[15:0]    reg_weight10_1_1;
wire[15:0]    reg_psum10_1_1;
wire[15:0]    reg_weight10_1_2;
wire[15:0]    reg_psum10_1_2;
wire[15:0]    reg_weight10_2_1;
wire[15:0]    reg_psum10_2_1;
wire[15:0]    reg_weight10_2_2;
wire[15:0]    reg_psum10_2_2;
wire[15:0]    reg_weight10_3_1;
wire[15:0]    reg_psum10_3_1;
wire[15:0]    reg_weight10_3_2;
wire[15:0]    reg_psum10_3_2;
wire[15:0]    reg_weight10_4_1;
wire[15:0]    reg_psum10_4_1;
wire[15:0]    reg_weight10_4_2;
wire[15:0]    reg_psum10_4_2;
wire[15:0]    reg_weight10_5_1;
wire[15:0]    reg_psum10_5_1;
wire[15:0]    reg_weight10_5_2;
wire[15:0]    reg_psum10_5_2;
wire[15:0]    reg_weight10_6_1;
wire[15:0]    reg_psum10_6_1;
wire[15:0]    reg_weight10_6_2;
wire[15:0]    reg_psum10_6_2;
wire[15:0]    reg_weight10_7_1;
wire[15:0]    reg_psum10_7_1;
wire[15:0]    reg_weight10_7_2;
wire[15:0]    reg_psum10_7_2;
wire[15:0]    reg_weight10_8_1;
wire[15:0]    reg_psum10_8_1;
wire[15:0]    reg_weight10_8_2;
wire[15:0]    reg_psum10_8_2;
wire[15:0]    reg_weight10_9_1;
wire[15:0]    reg_psum10_9_1;
wire[15:0]    reg_weight10_9_2;
wire[15:0]    reg_psum10_9_2;
wire[15:0]    reg_weight10_10_1;
wire[15:0]    reg_psum10_10_1;
wire[15:0]    reg_weight10_10_2;
wire[15:0]    reg_psum10_10_2;
wire[15:0]    reg_weight10_11_1;
wire[15:0]    reg_psum10_11_1;
wire[15:0]    reg_weight10_11_2;
wire[15:0]    reg_psum10_11_2;
wire[15:0]    reg_weight10_12_1;
wire[15:0]    reg_psum10_12_1;
wire[15:0]    reg_weight10_12_2;
wire[15:0]    reg_psum10_12_2;
wire[15:0]    reg_weight10_13_1;
wire[15:0]    reg_psum10_13_1;
wire[15:0]    reg_weight10_13_2;
wire[15:0]    reg_psum10_13_2;
wire[15:0]    reg_weight10_14_1;
wire[15:0]    reg_psum10_14_1;
wire[15:0]    reg_weight10_14_2;
wire[15:0]    reg_psum10_14_2;
wire[15:0]    reg_weight10_15_1;
wire[15:0]    reg_psum10_15_1;
wire[15:0]    reg_weight10_15_2;
wire[15:0]    reg_psum10_15_2;
wire[15:0]    reg_weight10_16_1;
wire[15:0]    reg_psum10_16_1;
wire[15:0]    reg_weight10_16_2;
wire[15:0]    reg_psum10_16_2;
wire[15:0]    reg_weight10_17_1;
wire[15:0]    reg_psum10_17_1;
wire[15:0]    reg_weight10_17_2;
wire[15:0]    reg_psum10_17_2;
wire[15:0]    reg_weight10_18_1;
wire[15:0]    reg_psum10_18_1;
wire[15:0]    reg_weight10_18_2;
wire[15:0]    reg_psum10_18_2;
wire[15:0]    reg_weight10_19_1;
wire[15:0]    reg_psum10_19_1;
wire[15:0]    reg_weight10_19_2;
wire[15:0]    reg_psum10_19_2;
wire[15:0]    reg_weight10_20_1;
wire[15:0]    reg_psum10_20_1;
wire[15:0]    reg_weight10_20_2;
wire[15:0]    reg_psum10_20_2;
wire[15:0]    reg_weight10_21_1;
wire[15:0]    reg_psum10_21_1;
wire[15:0]    reg_weight10_21_2;
wire[15:0]    reg_psum10_21_2;
wire[15:0]    reg_weight10_22_1;
wire[15:0]    reg_psum10_22_1;
wire[15:0]    reg_weight10_22_2;
wire[15:0]    reg_psum10_22_2;
wire[15:0]    reg_weight10_23_1;
wire[15:0]    reg_psum10_23_1;
wire[15:0]    reg_weight10_23_2;
wire[15:0]    reg_psum10_23_2;
wire[15:0]    reg_weight10_24_1;
wire[15:0]    reg_psum10_24_1;
wire[15:0]    reg_weight10_24_2;
wire[15:0]    reg_psum10_24_2;
wire[15:0]    reg_weight10_25_1;
wire[15:0]    reg_psum10_25_1;
wire[15:0]    reg_weight10_25_2;
wire[15:0]    reg_psum10_25_2;
wire[15:0]    reg_weight10_26_1;
wire[15:0]    reg_psum10_26_1;
wire[15:0]    reg_weight10_26_2;
wire[15:0]    reg_psum10_26_2;
wire[15:0]    reg_weight10_27_1;
wire[15:0]    reg_psum10_27_1;
wire[15:0]    reg_weight10_27_2;
wire[15:0]    reg_psum10_27_2;
wire[15:0]    reg_weight10_28_1;
wire[15:0]    reg_psum10_28_1;
wire[15:0]    reg_weight10_28_2;
wire[15:0]    reg_psum10_28_2;
wire[15:0]    reg_weight10_29_1;
wire[15:0]    reg_psum10_29_1;
wire[15:0]    reg_weight10_29_2;
wire[15:0]    reg_psum10_29_2;
wire[15:0]    reg_weight10_30_1;
wire[15:0]    reg_psum10_30_1;
wire[15:0]    reg_weight10_30_2;
wire[15:0]    reg_psum10_30_2;
wire[15:0]    reg_weight10_31_1;
wire[15:0]    reg_psum10_31_1;
wire[15:0]    reg_weight10_31_2;
wire[15:0]    reg_psum10_31_2;
wire[15:0]    reg_weight10_32_1;
wire[15:0]    reg_psum10_32_1;
wire[15:0]    reg_weight10_32_2;
wire[15:0]    reg_psum10_32_2;
wire[15:0]    reg_weight11_1_1;
wire[15:0]    reg_psum11_1_1;
wire[15:0]    reg_weight11_1_2;
wire[15:0]    reg_psum11_1_2;
wire[15:0]    reg_weight11_2_1;
wire[15:0]    reg_psum11_2_1;
wire[15:0]    reg_weight11_2_2;
wire[15:0]    reg_psum11_2_2;
wire[15:0]    reg_weight11_3_1;
wire[15:0]    reg_psum11_3_1;
wire[15:0]    reg_weight11_3_2;
wire[15:0]    reg_psum11_3_2;
wire[15:0]    reg_weight11_4_1;
wire[15:0]    reg_psum11_4_1;
wire[15:0]    reg_weight11_4_2;
wire[15:0]    reg_psum11_4_2;
wire[15:0]    reg_weight11_5_1;
wire[15:0]    reg_psum11_5_1;
wire[15:0]    reg_weight11_5_2;
wire[15:0]    reg_psum11_5_2;
wire[15:0]    reg_weight11_6_1;
wire[15:0]    reg_psum11_6_1;
wire[15:0]    reg_weight11_6_2;
wire[15:0]    reg_psum11_6_2;
wire[15:0]    reg_weight11_7_1;
wire[15:0]    reg_psum11_7_1;
wire[15:0]    reg_weight11_7_2;
wire[15:0]    reg_psum11_7_2;
wire[15:0]    reg_weight11_8_1;
wire[15:0]    reg_psum11_8_1;
wire[15:0]    reg_weight11_8_2;
wire[15:0]    reg_psum11_8_2;
wire[15:0]    reg_weight11_9_1;
wire[15:0]    reg_psum11_9_1;
wire[15:0]    reg_weight11_9_2;
wire[15:0]    reg_psum11_9_2;
wire[15:0]    reg_weight11_10_1;
wire[15:0]    reg_psum11_10_1;
wire[15:0]    reg_weight11_10_2;
wire[15:0]    reg_psum11_10_2;
wire[15:0]    reg_weight11_11_1;
wire[15:0]    reg_psum11_11_1;
wire[15:0]    reg_weight11_11_2;
wire[15:0]    reg_psum11_11_2;
wire[15:0]    reg_weight11_12_1;
wire[15:0]    reg_psum11_12_1;
wire[15:0]    reg_weight11_12_2;
wire[15:0]    reg_psum11_12_2;
wire[15:0]    reg_weight11_13_1;
wire[15:0]    reg_psum11_13_1;
wire[15:0]    reg_weight11_13_2;
wire[15:0]    reg_psum11_13_2;
wire[15:0]    reg_weight11_14_1;
wire[15:0]    reg_psum11_14_1;
wire[15:0]    reg_weight11_14_2;
wire[15:0]    reg_psum11_14_2;
wire[15:0]    reg_weight11_15_1;
wire[15:0]    reg_psum11_15_1;
wire[15:0]    reg_weight11_15_2;
wire[15:0]    reg_psum11_15_2;
wire[15:0]    reg_weight11_16_1;
wire[15:0]    reg_psum11_16_1;
wire[15:0]    reg_weight11_16_2;
wire[15:0]    reg_psum11_16_2;
wire[15:0]    reg_weight11_17_1;
wire[15:0]    reg_psum11_17_1;
wire[15:0]    reg_weight11_17_2;
wire[15:0]    reg_psum11_17_2;
wire[15:0]    reg_weight11_18_1;
wire[15:0]    reg_psum11_18_1;
wire[15:0]    reg_weight11_18_2;
wire[15:0]    reg_psum11_18_2;
wire[15:0]    reg_weight11_19_1;
wire[15:0]    reg_psum11_19_1;
wire[15:0]    reg_weight11_19_2;
wire[15:0]    reg_psum11_19_2;
wire[15:0]    reg_weight11_20_1;
wire[15:0]    reg_psum11_20_1;
wire[15:0]    reg_weight11_20_2;
wire[15:0]    reg_psum11_20_2;
wire[15:0]    reg_weight11_21_1;
wire[15:0]    reg_psum11_21_1;
wire[15:0]    reg_weight11_21_2;
wire[15:0]    reg_psum11_21_2;
wire[15:0]    reg_weight11_22_1;
wire[15:0]    reg_psum11_22_1;
wire[15:0]    reg_weight11_22_2;
wire[15:0]    reg_psum11_22_2;
wire[15:0]    reg_weight11_23_1;
wire[15:0]    reg_psum11_23_1;
wire[15:0]    reg_weight11_23_2;
wire[15:0]    reg_psum11_23_2;
wire[15:0]    reg_weight11_24_1;
wire[15:0]    reg_psum11_24_1;
wire[15:0]    reg_weight11_24_2;
wire[15:0]    reg_psum11_24_2;
wire[15:0]    reg_weight11_25_1;
wire[15:0]    reg_psum11_25_1;
wire[15:0]    reg_weight11_25_2;
wire[15:0]    reg_psum11_25_2;
wire[15:0]    reg_weight11_26_1;
wire[15:0]    reg_psum11_26_1;
wire[15:0]    reg_weight11_26_2;
wire[15:0]    reg_psum11_26_2;
wire[15:0]    reg_weight11_27_1;
wire[15:0]    reg_psum11_27_1;
wire[15:0]    reg_weight11_27_2;
wire[15:0]    reg_psum11_27_2;
wire[15:0]    reg_weight11_28_1;
wire[15:0]    reg_psum11_28_1;
wire[15:0]    reg_weight11_28_2;
wire[15:0]    reg_psum11_28_2;
wire[15:0]    reg_weight11_29_1;
wire[15:0]    reg_psum11_29_1;
wire[15:0]    reg_weight11_29_2;
wire[15:0]    reg_psum11_29_2;
wire[15:0]    reg_weight11_30_1;
wire[15:0]    reg_psum11_30_1;
wire[15:0]    reg_weight11_30_2;
wire[15:0]    reg_psum11_30_2;
wire[15:0]    reg_weight11_31_1;
wire[15:0]    reg_psum11_31_1;
wire[15:0]    reg_weight11_31_2;
wire[15:0]    reg_psum11_31_2;
wire[15:0]    reg_weight11_32_1;
wire[15:0]    reg_psum11_32_1;
wire[15:0]    reg_weight11_32_2;
wire[15:0]    reg_psum11_32_2;
wire[15:0]    reg_weight12_1_1;
wire[15:0]    reg_psum12_1_1;
wire[15:0]    reg_weight12_1_2;
wire[15:0]    reg_psum12_1_2;
wire[15:0]    reg_weight12_2_1;
wire[15:0]    reg_psum12_2_1;
wire[15:0]    reg_weight12_2_2;
wire[15:0]    reg_psum12_2_2;
wire[15:0]    reg_weight12_3_1;
wire[15:0]    reg_psum12_3_1;
wire[15:0]    reg_weight12_3_2;
wire[15:0]    reg_psum12_3_2;
wire[15:0]    reg_weight12_4_1;
wire[15:0]    reg_psum12_4_1;
wire[15:0]    reg_weight12_4_2;
wire[15:0]    reg_psum12_4_2;
wire[15:0]    reg_weight12_5_1;
wire[15:0]    reg_psum12_5_1;
wire[15:0]    reg_weight12_5_2;
wire[15:0]    reg_psum12_5_2;
wire[15:0]    reg_weight12_6_1;
wire[15:0]    reg_psum12_6_1;
wire[15:0]    reg_weight12_6_2;
wire[15:0]    reg_psum12_6_2;
wire[15:0]    reg_weight12_7_1;
wire[15:0]    reg_psum12_7_1;
wire[15:0]    reg_weight12_7_2;
wire[15:0]    reg_psum12_7_2;
wire[15:0]    reg_weight12_8_1;
wire[15:0]    reg_psum12_8_1;
wire[15:0]    reg_weight12_8_2;
wire[15:0]    reg_psum12_8_2;
wire[15:0]    reg_weight12_9_1;
wire[15:0]    reg_psum12_9_1;
wire[15:0]    reg_weight12_9_2;
wire[15:0]    reg_psum12_9_2;
wire[15:0]    reg_weight12_10_1;
wire[15:0]    reg_psum12_10_1;
wire[15:0]    reg_weight12_10_2;
wire[15:0]    reg_psum12_10_2;
wire[15:0]    reg_weight12_11_1;
wire[15:0]    reg_psum12_11_1;
wire[15:0]    reg_weight12_11_2;
wire[15:0]    reg_psum12_11_2;
wire[15:0]    reg_weight12_12_1;
wire[15:0]    reg_psum12_12_1;
wire[15:0]    reg_weight12_12_2;
wire[15:0]    reg_psum12_12_2;
wire[15:0]    reg_weight12_13_1;
wire[15:0]    reg_psum12_13_1;
wire[15:0]    reg_weight12_13_2;
wire[15:0]    reg_psum12_13_2;
wire[15:0]    reg_weight12_14_1;
wire[15:0]    reg_psum12_14_1;
wire[15:0]    reg_weight12_14_2;
wire[15:0]    reg_psum12_14_2;
wire[15:0]    reg_weight12_15_1;
wire[15:0]    reg_psum12_15_1;
wire[15:0]    reg_weight12_15_2;
wire[15:0]    reg_psum12_15_2;
wire[15:0]    reg_weight12_16_1;
wire[15:0]    reg_psum12_16_1;
wire[15:0]    reg_weight12_16_2;
wire[15:0]    reg_psum12_16_2;
wire[15:0]    reg_weight12_17_1;
wire[15:0]    reg_psum12_17_1;
wire[15:0]    reg_weight12_17_2;
wire[15:0]    reg_psum12_17_2;
wire[15:0]    reg_weight12_18_1;
wire[15:0]    reg_psum12_18_1;
wire[15:0]    reg_weight12_18_2;
wire[15:0]    reg_psum12_18_2;
wire[15:0]    reg_weight12_19_1;
wire[15:0]    reg_psum12_19_1;
wire[15:0]    reg_weight12_19_2;
wire[15:0]    reg_psum12_19_2;
wire[15:0]    reg_weight12_20_1;
wire[15:0]    reg_psum12_20_1;
wire[15:0]    reg_weight12_20_2;
wire[15:0]    reg_psum12_20_2;
wire[15:0]    reg_weight12_21_1;
wire[15:0]    reg_psum12_21_1;
wire[15:0]    reg_weight12_21_2;
wire[15:0]    reg_psum12_21_2;
wire[15:0]    reg_weight12_22_1;
wire[15:0]    reg_psum12_22_1;
wire[15:0]    reg_weight12_22_2;
wire[15:0]    reg_psum12_22_2;
wire[15:0]    reg_weight12_23_1;
wire[15:0]    reg_psum12_23_1;
wire[15:0]    reg_weight12_23_2;
wire[15:0]    reg_psum12_23_2;
wire[15:0]    reg_weight12_24_1;
wire[15:0]    reg_psum12_24_1;
wire[15:0]    reg_weight12_24_2;
wire[15:0]    reg_psum12_24_2;
wire[15:0]    reg_weight12_25_1;
wire[15:0]    reg_psum12_25_1;
wire[15:0]    reg_weight12_25_2;
wire[15:0]    reg_psum12_25_2;
wire[15:0]    reg_weight12_26_1;
wire[15:0]    reg_psum12_26_1;
wire[15:0]    reg_weight12_26_2;
wire[15:0]    reg_psum12_26_2;
wire[15:0]    reg_weight12_27_1;
wire[15:0]    reg_psum12_27_1;
wire[15:0]    reg_weight12_27_2;
wire[15:0]    reg_psum12_27_2;
wire[15:0]    reg_weight12_28_1;
wire[15:0]    reg_psum12_28_1;
wire[15:0]    reg_weight12_28_2;
wire[15:0]    reg_psum12_28_2;
wire[15:0]    reg_weight12_29_1;
wire[15:0]    reg_psum12_29_1;
wire[15:0]    reg_weight12_29_2;
wire[15:0]    reg_psum12_29_2;
wire[15:0]    reg_weight12_30_1;
wire[15:0]    reg_psum12_30_1;
wire[15:0]    reg_weight12_30_2;
wire[15:0]    reg_psum12_30_2;
wire[15:0]    reg_weight12_31_1;
wire[15:0]    reg_psum12_31_1;
wire[15:0]    reg_weight12_31_2;
wire[15:0]    reg_psum12_31_2;
wire[15:0]    reg_weight12_32_1;
wire[15:0]    reg_psum12_32_1;
wire[15:0]    reg_weight12_32_2;
wire[15:0]    reg_psum12_32_2;
wire[15:0]    reg_weight13_1_1;
wire[15:0]    reg_psum13_1_1;
wire[15:0]    reg_weight13_1_2;
wire[15:0]    reg_psum13_1_2;
wire[15:0]    reg_weight13_2_1;
wire[15:0]    reg_psum13_2_1;
wire[15:0]    reg_weight13_2_2;
wire[15:0]    reg_psum13_2_2;
wire[15:0]    reg_weight13_3_1;
wire[15:0]    reg_psum13_3_1;
wire[15:0]    reg_weight13_3_2;
wire[15:0]    reg_psum13_3_2;
wire[15:0]    reg_weight13_4_1;
wire[15:0]    reg_psum13_4_1;
wire[15:0]    reg_weight13_4_2;
wire[15:0]    reg_psum13_4_2;
wire[15:0]    reg_weight13_5_1;
wire[15:0]    reg_psum13_5_1;
wire[15:0]    reg_weight13_5_2;
wire[15:0]    reg_psum13_5_2;
wire[15:0]    reg_weight13_6_1;
wire[15:0]    reg_psum13_6_1;
wire[15:0]    reg_weight13_6_2;
wire[15:0]    reg_psum13_6_2;
wire[15:0]    reg_weight13_7_1;
wire[15:0]    reg_psum13_7_1;
wire[15:0]    reg_weight13_7_2;
wire[15:0]    reg_psum13_7_2;
wire[15:0]    reg_weight13_8_1;
wire[15:0]    reg_psum13_8_1;
wire[15:0]    reg_weight13_8_2;
wire[15:0]    reg_psum13_8_2;
wire[15:0]    reg_weight13_9_1;
wire[15:0]    reg_psum13_9_1;
wire[15:0]    reg_weight13_9_2;
wire[15:0]    reg_psum13_9_2;
wire[15:0]    reg_weight13_10_1;
wire[15:0]    reg_psum13_10_1;
wire[15:0]    reg_weight13_10_2;
wire[15:0]    reg_psum13_10_2;
wire[15:0]    reg_weight13_11_1;
wire[15:0]    reg_psum13_11_1;
wire[15:0]    reg_weight13_11_2;
wire[15:0]    reg_psum13_11_2;
wire[15:0]    reg_weight13_12_1;
wire[15:0]    reg_psum13_12_1;
wire[15:0]    reg_weight13_12_2;
wire[15:0]    reg_psum13_12_2;
wire[15:0]    reg_weight13_13_1;
wire[15:0]    reg_psum13_13_1;
wire[15:0]    reg_weight13_13_2;
wire[15:0]    reg_psum13_13_2;
wire[15:0]    reg_weight13_14_1;
wire[15:0]    reg_psum13_14_1;
wire[15:0]    reg_weight13_14_2;
wire[15:0]    reg_psum13_14_2;
wire[15:0]    reg_weight13_15_1;
wire[15:0]    reg_psum13_15_1;
wire[15:0]    reg_weight13_15_2;
wire[15:0]    reg_psum13_15_2;
wire[15:0]    reg_weight13_16_1;
wire[15:0]    reg_psum13_16_1;
wire[15:0]    reg_weight13_16_2;
wire[15:0]    reg_psum13_16_2;
wire[15:0]    reg_weight13_17_1;
wire[15:0]    reg_psum13_17_1;
wire[15:0]    reg_weight13_17_2;
wire[15:0]    reg_psum13_17_2;
wire[15:0]    reg_weight13_18_1;
wire[15:0]    reg_psum13_18_1;
wire[15:0]    reg_weight13_18_2;
wire[15:0]    reg_psum13_18_2;
wire[15:0]    reg_weight13_19_1;
wire[15:0]    reg_psum13_19_1;
wire[15:0]    reg_weight13_19_2;
wire[15:0]    reg_psum13_19_2;
wire[15:0]    reg_weight13_20_1;
wire[15:0]    reg_psum13_20_1;
wire[15:0]    reg_weight13_20_2;
wire[15:0]    reg_psum13_20_2;
wire[15:0]    reg_weight13_21_1;
wire[15:0]    reg_psum13_21_1;
wire[15:0]    reg_weight13_21_2;
wire[15:0]    reg_psum13_21_2;
wire[15:0]    reg_weight13_22_1;
wire[15:0]    reg_psum13_22_1;
wire[15:0]    reg_weight13_22_2;
wire[15:0]    reg_psum13_22_2;
wire[15:0]    reg_weight13_23_1;
wire[15:0]    reg_psum13_23_1;
wire[15:0]    reg_weight13_23_2;
wire[15:0]    reg_psum13_23_2;
wire[15:0]    reg_weight13_24_1;
wire[15:0]    reg_psum13_24_1;
wire[15:0]    reg_weight13_24_2;
wire[15:0]    reg_psum13_24_2;
wire[15:0]    reg_weight13_25_1;
wire[15:0]    reg_psum13_25_1;
wire[15:0]    reg_weight13_25_2;
wire[15:0]    reg_psum13_25_2;
wire[15:0]    reg_weight13_26_1;
wire[15:0]    reg_psum13_26_1;
wire[15:0]    reg_weight13_26_2;
wire[15:0]    reg_psum13_26_2;
wire[15:0]    reg_weight13_27_1;
wire[15:0]    reg_psum13_27_1;
wire[15:0]    reg_weight13_27_2;
wire[15:0]    reg_psum13_27_2;
wire[15:0]    reg_weight13_28_1;
wire[15:0]    reg_psum13_28_1;
wire[15:0]    reg_weight13_28_2;
wire[15:0]    reg_psum13_28_2;
wire[15:0]    reg_weight13_29_1;
wire[15:0]    reg_psum13_29_1;
wire[15:0]    reg_weight13_29_2;
wire[15:0]    reg_psum13_29_2;
wire[15:0]    reg_weight13_30_1;
wire[15:0]    reg_psum13_30_1;
wire[15:0]    reg_weight13_30_2;
wire[15:0]    reg_psum13_30_2;
wire[15:0]    reg_weight13_31_1;
wire[15:0]    reg_psum13_31_1;
wire[15:0]    reg_weight13_31_2;
wire[15:0]    reg_psum13_31_2;
wire[15:0]    reg_weight13_32_1;
wire[15:0]    reg_psum13_32_1;
wire[15:0]    reg_weight13_32_2;
wire[15:0]    reg_psum13_32_2;
wire[15:0]    reg_weight14_1_1;
wire[15:0]    reg_psum14_1_1;
wire[15:0]    reg_weight14_1_2;
wire[15:0]    reg_psum14_1_2;
wire[15:0]    reg_weight14_2_1;
wire[15:0]    reg_psum14_2_1;
wire[15:0]    reg_weight14_2_2;
wire[15:0]    reg_psum14_2_2;
wire[15:0]    reg_weight14_3_1;
wire[15:0]    reg_psum14_3_1;
wire[15:0]    reg_weight14_3_2;
wire[15:0]    reg_psum14_3_2;
wire[15:0]    reg_weight14_4_1;
wire[15:0]    reg_psum14_4_1;
wire[15:0]    reg_weight14_4_2;
wire[15:0]    reg_psum14_4_2;
wire[15:0]    reg_weight14_5_1;
wire[15:0]    reg_psum14_5_1;
wire[15:0]    reg_weight14_5_2;
wire[15:0]    reg_psum14_5_2;
wire[15:0]    reg_weight14_6_1;
wire[15:0]    reg_psum14_6_1;
wire[15:0]    reg_weight14_6_2;
wire[15:0]    reg_psum14_6_2;
wire[15:0]    reg_weight14_7_1;
wire[15:0]    reg_psum14_7_1;
wire[15:0]    reg_weight14_7_2;
wire[15:0]    reg_psum14_7_2;
wire[15:0]    reg_weight14_8_1;
wire[15:0]    reg_psum14_8_1;
wire[15:0]    reg_weight14_8_2;
wire[15:0]    reg_psum14_8_2;
wire[15:0]    reg_weight14_9_1;
wire[15:0]    reg_psum14_9_1;
wire[15:0]    reg_weight14_9_2;
wire[15:0]    reg_psum14_9_2;
wire[15:0]    reg_weight14_10_1;
wire[15:0]    reg_psum14_10_1;
wire[15:0]    reg_weight14_10_2;
wire[15:0]    reg_psum14_10_2;
wire[15:0]    reg_weight14_11_1;
wire[15:0]    reg_psum14_11_1;
wire[15:0]    reg_weight14_11_2;
wire[15:0]    reg_psum14_11_2;
wire[15:0]    reg_weight14_12_1;
wire[15:0]    reg_psum14_12_1;
wire[15:0]    reg_weight14_12_2;
wire[15:0]    reg_psum14_12_2;
wire[15:0]    reg_weight14_13_1;
wire[15:0]    reg_psum14_13_1;
wire[15:0]    reg_weight14_13_2;
wire[15:0]    reg_psum14_13_2;
wire[15:0]    reg_weight14_14_1;
wire[15:0]    reg_psum14_14_1;
wire[15:0]    reg_weight14_14_2;
wire[15:0]    reg_psum14_14_2;
wire[15:0]    reg_weight14_15_1;
wire[15:0]    reg_psum14_15_1;
wire[15:0]    reg_weight14_15_2;
wire[15:0]    reg_psum14_15_2;
wire[15:0]    reg_weight14_16_1;
wire[15:0]    reg_psum14_16_1;
wire[15:0]    reg_weight14_16_2;
wire[15:0]    reg_psum14_16_2;
wire[15:0]    reg_weight14_17_1;
wire[15:0]    reg_psum14_17_1;
wire[15:0]    reg_weight14_17_2;
wire[15:0]    reg_psum14_17_2;
wire[15:0]    reg_weight14_18_1;
wire[15:0]    reg_psum14_18_1;
wire[15:0]    reg_weight14_18_2;
wire[15:0]    reg_psum14_18_2;
wire[15:0]    reg_weight14_19_1;
wire[15:0]    reg_psum14_19_1;
wire[15:0]    reg_weight14_19_2;
wire[15:0]    reg_psum14_19_2;
wire[15:0]    reg_weight14_20_1;
wire[15:0]    reg_psum14_20_1;
wire[15:0]    reg_weight14_20_2;
wire[15:0]    reg_psum14_20_2;
wire[15:0]    reg_weight14_21_1;
wire[15:0]    reg_psum14_21_1;
wire[15:0]    reg_weight14_21_2;
wire[15:0]    reg_psum14_21_2;
wire[15:0]    reg_weight14_22_1;
wire[15:0]    reg_psum14_22_1;
wire[15:0]    reg_weight14_22_2;
wire[15:0]    reg_psum14_22_2;
wire[15:0]    reg_weight14_23_1;
wire[15:0]    reg_psum14_23_1;
wire[15:0]    reg_weight14_23_2;
wire[15:0]    reg_psum14_23_2;
wire[15:0]    reg_weight14_24_1;
wire[15:0]    reg_psum14_24_1;
wire[15:0]    reg_weight14_24_2;
wire[15:0]    reg_psum14_24_2;
wire[15:0]    reg_weight14_25_1;
wire[15:0]    reg_psum14_25_1;
wire[15:0]    reg_weight14_25_2;
wire[15:0]    reg_psum14_25_2;
wire[15:0]    reg_weight14_26_1;
wire[15:0]    reg_psum14_26_1;
wire[15:0]    reg_weight14_26_2;
wire[15:0]    reg_psum14_26_2;
wire[15:0]    reg_weight14_27_1;
wire[15:0]    reg_psum14_27_1;
wire[15:0]    reg_weight14_27_2;
wire[15:0]    reg_psum14_27_2;
wire[15:0]    reg_weight14_28_1;
wire[15:0]    reg_psum14_28_1;
wire[15:0]    reg_weight14_28_2;
wire[15:0]    reg_psum14_28_2;
wire[15:0]    reg_weight14_29_1;
wire[15:0]    reg_psum14_29_1;
wire[15:0]    reg_weight14_29_2;
wire[15:0]    reg_psum14_29_2;
wire[15:0]    reg_weight14_30_1;
wire[15:0]    reg_psum14_30_1;
wire[15:0]    reg_weight14_30_2;
wire[15:0]    reg_psum14_30_2;
wire[15:0]    reg_weight14_31_1;
wire[15:0]    reg_psum14_31_1;
wire[15:0]    reg_weight14_31_2;
wire[15:0]    reg_psum14_31_2;
wire[15:0]    reg_weight14_32_1;
wire[15:0]    reg_psum14_32_1;
wire[15:0]    reg_weight14_32_2;
wire[15:0]    reg_psum14_32_2;
wire[15:0]    reg_weight15_1_1;
wire[15:0]    reg_psum15_1_1;
wire[15:0]    reg_weight15_1_2;
wire[15:0]    reg_psum15_1_2;
wire[15:0]    reg_weight15_2_1;
wire[15:0]    reg_psum15_2_1;
wire[15:0]    reg_weight15_2_2;
wire[15:0]    reg_psum15_2_2;
wire[15:0]    reg_weight15_3_1;
wire[15:0]    reg_psum15_3_1;
wire[15:0]    reg_weight15_3_2;
wire[15:0]    reg_psum15_3_2;
wire[15:0]    reg_weight15_4_1;
wire[15:0]    reg_psum15_4_1;
wire[15:0]    reg_weight15_4_2;
wire[15:0]    reg_psum15_4_2;
wire[15:0]    reg_weight15_5_1;
wire[15:0]    reg_psum15_5_1;
wire[15:0]    reg_weight15_5_2;
wire[15:0]    reg_psum15_5_2;
wire[15:0]    reg_weight15_6_1;
wire[15:0]    reg_psum15_6_1;
wire[15:0]    reg_weight15_6_2;
wire[15:0]    reg_psum15_6_2;
wire[15:0]    reg_weight15_7_1;
wire[15:0]    reg_psum15_7_1;
wire[15:0]    reg_weight15_7_2;
wire[15:0]    reg_psum15_7_2;
wire[15:0]    reg_weight15_8_1;
wire[15:0]    reg_psum15_8_1;
wire[15:0]    reg_weight15_8_2;
wire[15:0]    reg_psum15_8_2;
wire[15:0]    reg_weight15_9_1;
wire[15:0]    reg_psum15_9_1;
wire[15:0]    reg_weight15_9_2;
wire[15:0]    reg_psum15_9_2;
wire[15:0]    reg_weight15_10_1;
wire[15:0]    reg_psum15_10_1;
wire[15:0]    reg_weight15_10_2;
wire[15:0]    reg_psum15_10_2;
wire[15:0]    reg_weight15_11_1;
wire[15:0]    reg_psum15_11_1;
wire[15:0]    reg_weight15_11_2;
wire[15:0]    reg_psum15_11_2;
wire[15:0]    reg_weight15_12_1;
wire[15:0]    reg_psum15_12_1;
wire[15:0]    reg_weight15_12_2;
wire[15:0]    reg_psum15_12_2;
wire[15:0]    reg_weight15_13_1;
wire[15:0]    reg_psum15_13_1;
wire[15:0]    reg_weight15_13_2;
wire[15:0]    reg_psum15_13_2;
wire[15:0]    reg_weight15_14_1;
wire[15:0]    reg_psum15_14_1;
wire[15:0]    reg_weight15_14_2;
wire[15:0]    reg_psum15_14_2;
wire[15:0]    reg_weight15_15_1;
wire[15:0]    reg_psum15_15_1;
wire[15:0]    reg_weight15_15_2;
wire[15:0]    reg_psum15_15_2;
wire[15:0]    reg_weight15_16_1;
wire[15:0]    reg_psum15_16_1;
wire[15:0]    reg_weight15_16_2;
wire[15:0]    reg_psum15_16_2;
wire[15:0]    reg_weight15_17_1;
wire[15:0]    reg_psum15_17_1;
wire[15:0]    reg_weight15_17_2;
wire[15:0]    reg_psum15_17_2;
wire[15:0]    reg_weight15_18_1;
wire[15:0]    reg_psum15_18_1;
wire[15:0]    reg_weight15_18_2;
wire[15:0]    reg_psum15_18_2;
wire[15:0]    reg_weight15_19_1;
wire[15:0]    reg_psum15_19_1;
wire[15:0]    reg_weight15_19_2;
wire[15:0]    reg_psum15_19_2;
wire[15:0]    reg_weight15_20_1;
wire[15:0]    reg_psum15_20_1;
wire[15:0]    reg_weight15_20_2;
wire[15:0]    reg_psum15_20_2;
wire[15:0]    reg_weight15_21_1;
wire[15:0]    reg_psum15_21_1;
wire[15:0]    reg_weight15_21_2;
wire[15:0]    reg_psum15_21_2;
wire[15:0]    reg_weight15_22_1;
wire[15:0]    reg_psum15_22_1;
wire[15:0]    reg_weight15_22_2;
wire[15:0]    reg_psum15_22_2;
wire[15:0]    reg_weight15_23_1;
wire[15:0]    reg_psum15_23_1;
wire[15:0]    reg_weight15_23_2;
wire[15:0]    reg_psum15_23_2;
wire[15:0]    reg_weight15_24_1;
wire[15:0]    reg_psum15_24_1;
wire[15:0]    reg_weight15_24_2;
wire[15:0]    reg_psum15_24_2;
wire[15:0]    reg_weight15_25_1;
wire[15:0]    reg_psum15_25_1;
wire[15:0]    reg_weight15_25_2;
wire[15:0]    reg_psum15_25_2;
wire[15:0]    reg_weight15_26_1;
wire[15:0]    reg_psum15_26_1;
wire[15:0]    reg_weight15_26_2;
wire[15:0]    reg_psum15_26_2;
wire[15:0]    reg_weight15_27_1;
wire[15:0]    reg_psum15_27_1;
wire[15:0]    reg_weight15_27_2;
wire[15:0]    reg_psum15_27_2;
wire[15:0]    reg_weight15_28_1;
wire[15:0]    reg_psum15_28_1;
wire[15:0]    reg_weight15_28_2;
wire[15:0]    reg_psum15_28_2;
wire[15:0]    reg_weight15_29_1;
wire[15:0]    reg_psum15_29_1;
wire[15:0]    reg_weight15_29_2;
wire[15:0]    reg_psum15_29_2;
wire[15:0]    reg_weight15_30_1;
wire[15:0]    reg_psum15_30_1;
wire[15:0]    reg_weight15_30_2;
wire[15:0]    reg_psum15_30_2;
wire[15:0]    reg_weight15_31_1;
wire[15:0]    reg_psum15_31_1;
wire[15:0]    reg_weight15_31_2;
wire[15:0]    reg_psum15_31_2;
wire[15:0]    reg_weight15_32_1;
wire[15:0]    reg_psum15_32_1;
wire[15:0]    reg_weight15_32_2;
wire[15:0]    reg_psum15_32_2;
wire[15:0]    reg_weight16_1_1;
wire[15:0]    reg_psum16_1_1;
wire[15:0]    reg_weight16_1_2;
wire[15:0]    reg_psum16_1_2;
wire[15:0]    reg_weight16_2_1;
wire[15:0]    reg_psum16_2_1;
wire[15:0]    reg_weight16_2_2;
wire[15:0]    reg_psum16_2_2;
wire[15:0]    reg_weight16_3_1;
wire[15:0]    reg_psum16_3_1;
wire[15:0]    reg_weight16_3_2;
wire[15:0]    reg_psum16_3_2;
wire[15:0]    reg_weight16_4_1;
wire[15:0]    reg_psum16_4_1;
wire[15:0]    reg_weight16_4_2;
wire[15:0]    reg_psum16_4_2;
wire[15:0]    reg_weight16_5_1;
wire[15:0]    reg_psum16_5_1;
wire[15:0]    reg_weight16_5_2;
wire[15:0]    reg_psum16_5_2;
wire[15:0]    reg_weight16_6_1;
wire[15:0]    reg_psum16_6_1;
wire[15:0]    reg_weight16_6_2;
wire[15:0]    reg_psum16_6_2;
wire[15:0]    reg_weight16_7_1;
wire[15:0]    reg_psum16_7_1;
wire[15:0]    reg_weight16_7_2;
wire[15:0]    reg_psum16_7_2;
wire[15:0]    reg_weight16_8_1;
wire[15:0]    reg_psum16_8_1;
wire[15:0]    reg_weight16_8_2;
wire[15:0]    reg_psum16_8_2;
wire[15:0]    reg_weight16_9_1;
wire[15:0]    reg_psum16_9_1;
wire[15:0]    reg_weight16_9_2;
wire[15:0]    reg_psum16_9_2;
wire[15:0]    reg_weight16_10_1;
wire[15:0]    reg_psum16_10_1;
wire[15:0]    reg_weight16_10_2;
wire[15:0]    reg_psum16_10_2;
wire[15:0]    reg_weight16_11_1;
wire[15:0]    reg_psum16_11_1;
wire[15:0]    reg_weight16_11_2;
wire[15:0]    reg_psum16_11_2;
wire[15:0]    reg_weight16_12_1;
wire[15:0]    reg_psum16_12_1;
wire[15:0]    reg_weight16_12_2;
wire[15:0]    reg_psum16_12_2;
wire[15:0]    reg_weight16_13_1;
wire[15:0]    reg_psum16_13_1;
wire[15:0]    reg_weight16_13_2;
wire[15:0]    reg_psum16_13_2;
wire[15:0]    reg_weight16_14_1;
wire[15:0]    reg_psum16_14_1;
wire[15:0]    reg_weight16_14_2;
wire[15:0]    reg_psum16_14_2;
wire[15:0]    reg_weight16_15_1;
wire[15:0]    reg_psum16_15_1;
wire[15:0]    reg_weight16_15_2;
wire[15:0]    reg_psum16_15_2;
wire[15:0]    reg_weight16_16_1;
wire[15:0]    reg_psum16_16_1;
wire[15:0]    reg_weight16_16_2;
wire[15:0]    reg_psum16_16_2;
wire[15:0]    reg_weight16_17_1;
wire[15:0]    reg_psum16_17_1;
wire[15:0]    reg_weight16_17_2;
wire[15:0]    reg_psum16_17_2;
wire[15:0]    reg_weight16_18_1;
wire[15:0]    reg_psum16_18_1;
wire[15:0]    reg_weight16_18_2;
wire[15:0]    reg_psum16_18_2;
wire[15:0]    reg_weight16_19_1;
wire[15:0]    reg_psum16_19_1;
wire[15:0]    reg_weight16_19_2;
wire[15:0]    reg_psum16_19_2;
wire[15:0]    reg_weight16_20_1;
wire[15:0]    reg_psum16_20_1;
wire[15:0]    reg_weight16_20_2;
wire[15:0]    reg_psum16_20_2;
wire[15:0]    reg_weight16_21_1;
wire[15:0]    reg_psum16_21_1;
wire[15:0]    reg_weight16_21_2;
wire[15:0]    reg_psum16_21_2;
wire[15:0]    reg_weight16_22_1;
wire[15:0]    reg_psum16_22_1;
wire[15:0]    reg_weight16_22_2;
wire[15:0]    reg_psum16_22_2;
wire[15:0]    reg_weight16_23_1;
wire[15:0]    reg_psum16_23_1;
wire[15:0]    reg_weight16_23_2;
wire[15:0]    reg_psum16_23_2;
wire[15:0]    reg_weight16_24_1;
wire[15:0]    reg_psum16_24_1;
wire[15:0]    reg_weight16_24_2;
wire[15:0]    reg_psum16_24_2;
wire[15:0]    reg_weight16_25_1;
wire[15:0]    reg_psum16_25_1;
wire[15:0]    reg_weight16_25_2;
wire[15:0]    reg_psum16_25_2;
wire[15:0]    reg_weight16_26_1;
wire[15:0]    reg_psum16_26_1;
wire[15:0]    reg_weight16_26_2;
wire[15:0]    reg_psum16_26_2;
wire[15:0]    reg_weight16_27_1;
wire[15:0]    reg_psum16_27_1;
wire[15:0]    reg_weight16_27_2;
wire[15:0]    reg_psum16_27_2;
wire[15:0]    reg_weight16_28_1;
wire[15:0]    reg_psum16_28_1;
wire[15:0]    reg_weight16_28_2;
wire[15:0]    reg_psum16_28_2;
wire[15:0]    reg_weight16_29_1;
wire[15:0]    reg_psum16_29_1;
wire[15:0]    reg_weight16_29_2;
wire[15:0]    reg_psum16_29_2;
wire[15:0]    reg_weight16_30_1;
wire[15:0]    reg_psum16_30_1;
wire[15:0]    reg_weight16_30_2;
wire[15:0]    reg_psum16_30_2;
wire[15:0]    reg_weight16_31_1;
wire[15:0]    reg_psum16_31_1;
wire[15:0]    reg_weight16_31_2;
wire[15:0]    reg_psum16_31_2;
wire[15:0]    reg_weight16_32_1;
wire[15:0]    reg_psum16_32_1;
wire[15:0]    reg_weight16_32_2;
wire[15:0]    reg_psum16_32_2;
wire[15:0]    reg_weight17_1_1;
wire[15:0]    reg_psum17_1_1;
wire[15:0]    reg_weight17_1_2;
wire[15:0]    reg_psum17_1_2;
wire[15:0]    reg_weight17_2_1;
wire[15:0]    reg_psum17_2_1;
wire[15:0]    reg_weight17_2_2;
wire[15:0]    reg_psum17_2_2;
wire[15:0]    reg_weight17_3_1;
wire[15:0]    reg_psum17_3_1;
wire[15:0]    reg_weight17_3_2;
wire[15:0]    reg_psum17_3_2;
wire[15:0]    reg_weight17_4_1;
wire[15:0]    reg_psum17_4_1;
wire[15:0]    reg_weight17_4_2;
wire[15:0]    reg_psum17_4_2;
wire[15:0]    reg_weight17_5_1;
wire[15:0]    reg_psum17_5_1;
wire[15:0]    reg_weight17_5_2;
wire[15:0]    reg_psum17_5_2;
wire[15:0]    reg_weight17_6_1;
wire[15:0]    reg_psum17_6_1;
wire[15:0]    reg_weight17_6_2;
wire[15:0]    reg_psum17_6_2;
wire[15:0]    reg_weight17_7_1;
wire[15:0]    reg_psum17_7_1;
wire[15:0]    reg_weight17_7_2;
wire[15:0]    reg_psum17_7_2;
wire[15:0]    reg_weight17_8_1;
wire[15:0]    reg_psum17_8_1;
wire[15:0]    reg_weight17_8_2;
wire[15:0]    reg_psum17_8_2;
wire[15:0]    reg_weight17_9_1;
wire[15:0]    reg_psum17_9_1;
wire[15:0]    reg_weight17_9_2;
wire[15:0]    reg_psum17_9_2;
wire[15:0]    reg_weight17_10_1;
wire[15:0]    reg_psum17_10_1;
wire[15:0]    reg_weight17_10_2;
wire[15:0]    reg_psum17_10_2;
wire[15:0]    reg_weight17_11_1;
wire[15:0]    reg_psum17_11_1;
wire[15:0]    reg_weight17_11_2;
wire[15:0]    reg_psum17_11_2;
wire[15:0]    reg_weight17_12_1;
wire[15:0]    reg_psum17_12_1;
wire[15:0]    reg_weight17_12_2;
wire[15:0]    reg_psum17_12_2;
wire[15:0]    reg_weight17_13_1;
wire[15:0]    reg_psum17_13_1;
wire[15:0]    reg_weight17_13_2;
wire[15:0]    reg_psum17_13_2;
wire[15:0]    reg_weight17_14_1;
wire[15:0]    reg_psum17_14_1;
wire[15:0]    reg_weight17_14_2;
wire[15:0]    reg_psum17_14_2;
wire[15:0]    reg_weight17_15_1;
wire[15:0]    reg_psum17_15_1;
wire[15:0]    reg_weight17_15_2;
wire[15:0]    reg_psum17_15_2;
wire[15:0]    reg_weight17_16_1;
wire[15:0]    reg_psum17_16_1;
wire[15:0]    reg_weight17_16_2;
wire[15:0]    reg_psum17_16_2;
wire[15:0]    reg_weight17_17_1;
wire[15:0]    reg_psum17_17_1;
wire[15:0]    reg_weight17_17_2;
wire[15:0]    reg_psum17_17_2;
wire[15:0]    reg_weight17_18_1;
wire[15:0]    reg_psum17_18_1;
wire[15:0]    reg_weight17_18_2;
wire[15:0]    reg_psum17_18_2;
wire[15:0]    reg_weight17_19_1;
wire[15:0]    reg_psum17_19_1;
wire[15:0]    reg_weight17_19_2;
wire[15:0]    reg_psum17_19_2;
wire[15:0]    reg_weight17_20_1;
wire[15:0]    reg_psum17_20_1;
wire[15:0]    reg_weight17_20_2;
wire[15:0]    reg_psum17_20_2;
wire[15:0]    reg_weight17_21_1;
wire[15:0]    reg_psum17_21_1;
wire[15:0]    reg_weight17_21_2;
wire[15:0]    reg_psum17_21_2;
wire[15:0]    reg_weight17_22_1;
wire[15:0]    reg_psum17_22_1;
wire[15:0]    reg_weight17_22_2;
wire[15:0]    reg_psum17_22_2;
wire[15:0]    reg_weight17_23_1;
wire[15:0]    reg_psum17_23_1;
wire[15:0]    reg_weight17_23_2;
wire[15:0]    reg_psum17_23_2;
wire[15:0]    reg_weight17_24_1;
wire[15:0]    reg_psum17_24_1;
wire[15:0]    reg_weight17_24_2;
wire[15:0]    reg_psum17_24_2;
wire[15:0]    reg_weight17_25_1;
wire[15:0]    reg_psum17_25_1;
wire[15:0]    reg_weight17_25_2;
wire[15:0]    reg_psum17_25_2;
wire[15:0]    reg_weight17_26_1;
wire[15:0]    reg_psum17_26_1;
wire[15:0]    reg_weight17_26_2;
wire[15:0]    reg_psum17_26_2;
wire[15:0]    reg_weight17_27_1;
wire[15:0]    reg_psum17_27_1;
wire[15:0]    reg_weight17_27_2;
wire[15:0]    reg_psum17_27_2;
wire[15:0]    reg_weight17_28_1;
wire[15:0]    reg_psum17_28_1;
wire[15:0]    reg_weight17_28_2;
wire[15:0]    reg_psum17_28_2;
wire[15:0]    reg_weight17_29_1;
wire[15:0]    reg_psum17_29_1;
wire[15:0]    reg_weight17_29_2;
wire[15:0]    reg_psum17_29_2;
wire[15:0]    reg_weight17_30_1;
wire[15:0]    reg_psum17_30_1;
wire[15:0]    reg_weight17_30_2;
wire[15:0]    reg_psum17_30_2;
wire[15:0]    reg_weight17_31_1;
wire[15:0]    reg_psum17_31_1;
wire[15:0]    reg_weight17_31_2;
wire[15:0]    reg_psum17_31_2;
wire[15:0]    reg_weight17_32_1;
wire[15:0]    reg_psum17_32_1;
wire[15:0]    reg_weight17_32_2;
wire[15:0]    reg_psum17_32_2;
wire[15:0]    reg_weight18_1_1;
wire[15:0]    reg_psum18_1_1;
wire[15:0]    reg_weight18_1_2;
wire[15:0]    reg_psum18_1_2;
wire[15:0]    reg_weight18_2_1;
wire[15:0]    reg_psum18_2_1;
wire[15:0]    reg_weight18_2_2;
wire[15:0]    reg_psum18_2_2;
wire[15:0]    reg_weight18_3_1;
wire[15:0]    reg_psum18_3_1;
wire[15:0]    reg_weight18_3_2;
wire[15:0]    reg_psum18_3_2;
wire[15:0]    reg_weight18_4_1;
wire[15:0]    reg_psum18_4_1;
wire[15:0]    reg_weight18_4_2;
wire[15:0]    reg_psum18_4_2;
wire[15:0]    reg_weight18_5_1;
wire[15:0]    reg_psum18_5_1;
wire[15:0]    reg_weight18_5_2;
wire[15:0]    reg_psum18_5_2;
wire[15:0]    reg_weight18_6_1;
wire[15:0]    reg_psum18_6_1;
wire[15:0]    reg_weight18_6_2;
wire[15:0]    reg_psum18_6_2;
wire[15:0]    reg_weight18_7_1;
wire[15:0]    reg_psum18_7_1;
wire[15:0]    reg_weight18_7_2;
wire[15:0]    reg_psum18_7_2;
wire[15:0]    reg_weight18_8_1;
wire[15:0]    reg_psum18_8_1;
wire[15:0]    reg_weight18_8_2;
wire[15:0]    reg_psum18_8_2;
wire[15:0]    reg_weight18_9_1;
wire[15:0]    reg_psum18_9_1;
wire[15:0]    reg_weight18_9_2;
wire[15:0]    reg_psum18_9_2;
wire[15:0]    reg_weight18_10_1;
wire[15:0]    reg_psum18_10_1;
wire[15:0]    reg_weight18_10_2;
wire[15:0]    reg_psum18_10_2;
wire[15:0]    reg_weight18_11_1;
wire[15:0]    reg_psum18_11_1;
wire[15:0]    reg_weight18_11_2;
wire[15:0]    reg_psum18_11_2;
wire[15:0]    reg_weight18_12_1;
wire[15:0]    reg_psum18_12_1;
wire[15:0]    reg_weight18_12_2;
wire[15:0]    reg_psum18_12_2;
wire[15:0]    reg_weight18_13_1;
wire[15:0]    reg_psum18_13_1;
wire[15:0]    reg_weight18_13_2;
wire[15:0]    reg_psum18_13_2;
wire[15:0]    reg_weight18_14_1;
wire[15:0]    reg_psum18_14_1;
wire[15:0]    reg_weight18_14_2;
wire[15:0]    reg_psum18_14_2;
wire[15:0]    reg_weight18_15_1;
wire[15:0]    reg_psum18_15_1;
wire[15:0]    reg_weight18_15_2;
wire[15:0]    reg_psum18_15_2;
wire[15:0]    reg_weight18_16_1;
wire[15:0]    reg_psum18_16_1;
wire[15:0]    reg_weight18_16_2;
wire[15:0]    reg_psum18_16_2;
wire[15:0]    reg_weight18_17_1;
wire[15:0]    reg_psum18_17_1;
wire[15:0]    reg_weight18_17_2;
wire[15:0]    reg_psum18_17_2;
wire[15:0]    reg_weight18_18_1;
wire[15:0]    reg_psum18_18_1;
wire[15:0]    reg_weight18_18_2;
wire[15:0]    reg_psum18_18_2;
wire[15:0]    reg_weight18_19_1;
wire[15:0]    reg_psum18_19_1;
wire[15:0]    reg_weight18_19_2;
wire[15:0]    reg_psum18_19_2;
wire[15:0]    reg_weight18_20_1;
wire[15:0]    reg_psum18_20_1;
wire[15:0]    reg_weight18_20_2;
wire[15:0]    reg_psum18_20_2;
wire[15:0]    reg_weight18_21_1;
wire[15:0]    reg_psum18_21_1;
wire[15:0]    reg_weight18_21_2;
wire[15:0]    reg_psum18_21_2;
wire[15:0]    reg_weight18_22_1;
wire[15:0]    reg_psum18_22_1;
wire[15:0]    reg_weight18_22_2;
wire[15:0]    reg_psum18_22_2;
wire[15:0]    reg_weight18_23_1;
wire[15:0]    reg_psum18_23_1;
wire[15:0]    reg_weight18_23_2;
wire[15:0]    reg_psum18_23_2;
wire[15:0]    reg_weight18_24_1;
wire[15:0]    reg_psum18_24_1;
wire[15:0]    reg_weight18_24_2;
wire[15:0]    reg_psum18_24_2;
wire[15:0]    reg_weight18_25_1;
wire[15:0]    reg_psum18_25_1;
wire[15:0]    reg_weight18_25_2;
wire[15:0]    reg_psum18_25_2;
wire[15:0]    reg_weight18_26_1;
wire[15:0]    reg_psum18_26_1;
wire[15:0]    reg_weight18_26_2;
wire[15:0]    reg_psum18_26_2;
wire[15:0]    reg_weight18_27_1;
wire[15:0]    reg_psum18_27_1;
wire[15:0]    reg_weight18_27_2;
wire[15:0]    reg_psum18_27_2;
wire[15:0]    reg_weight18_28_1;
wire[15:0]    reg_psum18_28_1;
wire[15:0]    reg_weight18_28_2;
wire[15:0]    reg_psum18_28_2;
wire[15:0]    reg_weight18_29_1;
wire[15:0]    reg_psum18_29_1;
wire[15:0]    reg_weight18_29_2;
wire[15:0]    reg_psum18_29_2;
wire[15:0]    reg_weight18_30_1;
wire[15:0]    reg_psum18_30_1;
wire[15:0]    reg_weight18_30_2;
wire[15:0]    reg_psum18_30_2;
wire[15:0]    reg_weight18_31_1;
wire[15:0]    reg_psum18_31_1;
wire[15:0]    reg_weight18_31_2;
wire[15:0]    reg_psum18_31_2;
wire[15:0]    reg_weight18_32_1;
wire[15:0]    reg_psum18_32_1;
wire[15:0]    reg_weight18_32_2;
wire[15:0]    reg_psum18_32_2;
wire[15:0]    reg_weight19_1_1;
wire[15:0]    reg_psum19_1_1;
wire[15:0]    reg_weight19_1_2;
wire[15:0]    reg_psum19_1_2;
wire[15:0]    reg_weight19_2_1;
wire[15:0]    reg_psum19_2_1;
wire[15:0]    reg_weight19_2_2;
wire[15:0]    reg_psum19_2_2;
wire[15:0]    reg_weight19_3_1;
wire[15:0]    reg_psum19_3_1;
wire[15:0]    reg_weight19_3_2;
wire[15:0]    reg_psum19_3_2;
wire[15:0]    reg_weight19_4_1;
wire[15:0]    reg_psum19_4_1;
wire[15:0]    reg_weight19_4_2;
wire[15:0]    reg_psum19_4_2;
wire[15:0]    reg_weight19_5_1;
wire[15:0]    reg_psum19_5_1;
wire[15:0]    reg_weight19_5_2;
wire[15:0]    reg_psum19_5_2;
wire[15:0]    reg_weight19_6_1;
wire[15:0]    reg_psum19_6_1;
wire[15:0]    reg_weight19_6_2;
wire[15:0]    reg_psum19_6_2;
wire[15:0]    reg_weight19_7_1;
wire[15:0]    reg_psum19_7_1;
wire[15:0]    reg_weight19_7_2;
wire[15:0]    reg_psum19_7_2;
wire[15:0]    reg_weight19_8_1;
wire[15:0]    reg_psum19_8_1;
wire[15:0]    reg_weight19_8_2;
wire[15:0]    reg_psum19_8_2;
wire[15:0]    reg_weight19_9_1;
wire[15:0]    reg_psum19_9_1;
wire[15:0]    reg_weight19_9_2;
wire[15:0]    reg_psum19_9_2;
wire[15:0]    reg_weight19_10_1;
wire[15:0]    reg_psum19_10_1;
wire[15:0]    reg_weight19_10_2;
wire[15:0]    reg_psum19_10_2;
wire[15:0]    reg_weight19_11_1;
wire[15:0]    reg_psum19_11_1;
wire[15:0]    reg_weight19_11_2;
wire[15:0]    reg_psum19_11_2;
wire[15:0]    reg_weight19_12_1;
wire[15:0]    reg_psum19_12_1;
wire[15:0]    reg_weight19_12_2;
wire[15:0]    reg_psum19_12_2;
wire[15:0]    reg_weight19_13_1;
wire[15:0]    reg_psum19_13_1;
wire[15:0]    reg_weight19_13_2;
wire[15:0]    reg_psum19_13_2;
wire[15:0]    reg_weight19_14_1;
wire[15:0]    reg_psum19_14_1;
wire[15:0]    reg_weight19_14_2;
wire[15:0]    reg_psum19_14_2;
wire[15:0]    reg_weight19_15_1;
wire[15:0]    reg_psum19_15_1;
wire[15:0]    reg_weight19_15_2;
wire[15:0]    reg_psum19_15_2;
wire[15:0]    reg_weight19_16_1;
wire[15:0]    reg_psum19_16_1;
wire[15:0]    reg_weight19_16_2;
wire[15:0]    reg_psum19_16_2;
wire[15:0]    reg_weight19_17_1;
wire[15:0]    reg_psum19_17_1;
wire[15:0]    reg_weight19_17_2;
wire[15:0]    reg_psum19_17_2;
wire[15:0]    reg_weight19_18_1;
wire[15:0]    reg_psum19_18_1;
wire[15:0]    reg_weight19_18_2;
wire[15:0]    reg_psum19_18_2;
wire[15:0]    reg_weight19_19_1;
wire[15:0]    reg_psum19_19_1;
wire[15:0]    reg_weight19_19_2;
wire[15:0]    reg_psum19_19_2;
wire[15:0]    reg_weight19_20_1;
wire[15:0]    reg_psum19_20_1;
wire[15:0]    reg_weight19_20_2;
wire[15:0]    reg_psum19_20_2;
wire[15:0]    reg_weight19_21_1;
wire[15:0]    reg_psum19_21_1;
wire[15:0]    reg_weight19_21_2;
wire[15:0]    reg_psum19_21_2;
wire[15:0]    reg_weight19_22_1;
wire[15:0]    reg_psum19_22_1;
wire[15:0]    reg_weight19_22_2;
wire[15:0]    reg_psum19_22_2;
wire[15:0]    reg_weight19_23_1;
wire[15:0]    reg_psum19_23_1;
wire[15:0]    reg_weight19_23_2;
wire[15:0]    reg_psum19_23_2;
wire[15:0]    reg_weight19_24_1;
wire[15:0]    reg_psum19_24_1;
wire[15:0]    reg_weight19_24_2;
wire[15:0]    reg_psum19_24_2;
wire[15:0]    reg_weight19_25_1;
wire[15:0]    reg_psum19_25_1;
wire[15:0]    reg_weight19_25_2;
wire[15:0]    reg_psum19_25_2;
wire[15:0]    reg_weight19_26_1;
wire[15:0]    reg_psum19_26_1;
wire[15:0]    reg_weight19_26_2;
wire[15:0]    reg_psum19_26_2;
wire[15:0]    reg_weight19_27_1;
wire[15:0]    reg_psum19_27_1;
wire[15:0]    reg_weight19_27_2;
wire[15:0]    reg_psum19_27_2;
wire[15:0]    reg_weight19_28_1;
wire[15:0]    reg_psum19_28_1;
wire[15:0]    reg_weight19_28_2;
wire[15:0]    reg_psum19_28_2;
wire[15:0]    reg_weight19_29_1;
wire[15:0]    reg_psum19_29_1;
wire[15:0]    reg_weight19_29_2;
wire[15:0]    reg_psum19_29_2;
wire[15:0]    reg_weight19_30_1;
wire[15:0]    reg_psum19_30_1;
wire[15:0]    reg_weight19_30_2;
wire[15:0]    reg_psum19_30_2;
wire[15:0]    reg_weight19_31_1;
wire[15:0]    reg_psum19_31_1;
wire[15:0]    reg_weight19_31_2;
wire[15:0]    reg_psum19_31_2;
wire[15:0]    reg_weight19_32_1;
wire[15:0]    reg_psum19_32_1;
wire[15:0]    reg_weight19_32_2;
wire[15:0]    reg_psum19_32_2;
wire[15:0]    reg_weight20_1_1;
wire[15:0]    reg_psum20_1_1;
wire[15:0]    reg_weight20_1_2;
wire[15:0]    reg_psum20_1_2;
wire[15:0]    reg_weight20_2_1;
wire[15:0]    reg_psum20_2_1;
wire[15:0]    reg_weight20_2_2;
wire[15:0]    reg_psum20_2_2;
wire[15:0]    reg_weight20_3_1;
wire[15:0]    reg_psum20_3_1;
wire[15:0]    reg_weight20_3_2;
wire[15:0]    reg_psum20_3_2;
wire[15:0]    reg_weight20_4_1;
wire[15:0]    reg_psum20_4_1;
wire[15:0]    reg_weight20_4_2;
wire[15:0]    reg_psum20_4_2;
wire[15:0]    reg_weight20_5_1;
wire[15:0]    reg_psum20_5_1;
wire[15:0]    reg_weight20_5_2;
wire[15:0]    reg_psum20_5_2;
wire[15:0]    reg_weight20_6_1;
wire[15:0]    reg_psum20_6_1;
wire[15:0]    reg_weight20_6_2;
wire[15:0]    reg_psum20_6_2;
wire[15:0]    reg_weight20_7_1;
wire[15:0]    reg_psum20_7_1;
wire[15:0]    reg_weight20_7_2;
wire[15:0]    reg_psum20_7_2;
wire[15:0]    reg_weight20_8_1;
wire[15:0]    reg_psum20_8_1;
wire[15:0]    reg_weight20_8_2;
wire[15:0]    reg_psum20_8_2;
wire[15:0]    reg_weight20_9_1;
wire[15:0]    reg_psum20_9_1;
wire[15:0]    reg_weight20_9_2;
wire[15:0]    reg_psum20_9_2;
wire[15:0]    reg_weight20_10_1;
wire[15:0]    reg_psum20_10_1;
wire[15:0]    reg_weight20_10_2;
wire[15:0]    reg_psum20_10_2;
wire[15:0]    reg_weight20_11_1;
wire[15:0]    reg_psum20_11_1;
wire[15:0]    reg_weight20_11_2;
wire[15:0]    reg_psum20_11_2;
wire[15:0]    reg_weight20_12_1;
wire[15:0]    reg_psum20_12_1;
wire[15:0]    reg_weight20_12_2;
wire[15:0]    reg_psum20_12_2;
wire[15:0]    reg_weight20_13_1;
wire[15:0]    reg_psum20_13_1;
wire[15:0]    reg_weight20_13_2;
wire[15:0]    reg_psum20_13_2;
wire[15:0]    reg_weight20_14_1;
wire[15:0]    reg_psum20_14_1;
wire[15:0]    reg_weight20_14_2;
wire[15:0]    reg_psum20_14_2;
wire[15:0]    reg_weight20_15_1;
wire[15:0]    reg_psum20_15_1;
wire[15:0]    reg_weight20_15_2;
wire[15:0]    reg_psum20_15_2;
wire[15:0]    reg_weight20_16_1;
wire[15:0]    reg_psum20_16_1;
wire[15:0]    reg_weight20_16_2;
wire[15:0]    reg_psum20_16_2;
wire[15:0]    reg_weight20_17_1;
wire[15:0]    reg_psum20_17_1;
wire[15:0]    reg_weight20_17_2;
wire[15:0]    reg_psum20_17_2;
wire[15:0]    reg_weight20_18_1;
wire[15:0]    reg_psum20_18_1;
wire[15:0]    reg_weight20_18_2;
wire[15:0]    reg_psum20_18_2;
wire[15:0]    reg_weight20_19_1;
wire[15:0]    reg_psum20_19_1;
wire[15:0]    reg_weight20_19_2;
wire[15:0]    reg_psum20_19_2;
wire[15:0]    reg_weight20_20_1;
wire[15:0]    reg_psum20_20_1;
wire[15:0]    reg_weight20_20_2;
wire[15:0]    reg_psum20_20_2;
wire[15:0]    reg_weight20_21_1;
wire[15:0]    reg_psum20_21_1;
wire[15:0]    reg_weight20_21_2;
wire[15:0]    reg_psum20_21_2;
wire[15:0]    reg_weight20_22_1;
wire[15:0]    reg_psum20_22_1;
wire[15:0]    reg_weight20_22_2;
wire[15:0]    reg_psum20_22_2;
wire[15:0]    reg_weight20_23_1;
wire[15:0]    reg_psum20_23_1;
wire[15:0]    reg_weight20_23_2;
wire[15:0]    reg_psum20_23_2;
wire[15:0]    reg_weight20_24_1;
wire[15:0]    reg_psum20_24_1;
wire[15:0]    reg_weight20_24_2;
wire[15:0]    reg_psum20_24_2;
wire[15:0]    reg_weight20_25_1;
wire[15:0]    reg_psum20_25_1;
wire[15:0]    reg_weight20_25_2;
wire[15:0]    reg_psum20_25_2;
wire[15:0]    reg_weight20_26_1;
wire[15:0]    reg_psum20_26_1;
wire[15:0]    reg_weight20_26_2;
wire[15:0]    reg_psum20_26_2;
wire[15:0]    reg_weight20_27_1;
wire[15:0]    reg_psum20_27_1;
wire[15:0]    reg_weight20_27_2;
wire[15:0]    reg_psum20_27_2;
wire[15:0]    reg_weight20_28_1;
wire[15:0]    reg_psum20_28_1;
wire[15:0]    reg_weight20_28_2;
wire[15:0]    reg_psum20_28_2;
wire[15:0]    reg_weight20_29_1;
wire[15:0]    reg_psum20_29_1;
wire[15:0]    reg_weight20_29_2;
wire[15:0]    reg_psum20_29_2;
wire[15:0]    reg_weight20_30_1;
wire[15:0]    reg_psum20_30_1;
wire[15:0]    reg_weight20_30_2;
wire[15:0]    reg_psum20_30_2;
wire[15:0]    reg_weight20_31_1;
wire[15:0]    reg_psum20_31_1;
wire[15:0]    reg_weight20_31_2;
wire[15:0]    reg_psum20_31_2;
wire[15:0]    reg_weight20_32_1;
wire[15:0]    reg_psum20_32_1;
wire[15:0]    reg_weight20_32_2;
wire[15:0]    reg_psum20_32_2;
wire[15:0]    reg_weight21_1_1;
wire[15:0]    reg_psum21_1_1;
wire[15:0]    reg_weight21_1_2;
wire[15:0]    reg_psum21_1_2;
wire[15:0]    reg_weight21_2_1;
wire[15:0]    reg_psum21_2_1;
wire[15:0]    reg_weight21_2_2;
wire[15:0]    reg_psum21_2_2;
wire[15:0]    reg_weight21_3_1;
wire[15:0]    reg_psum21_3_1;
wire[15:0]    reg_weight21_3_2;
wire[15:0]    reg_psum21_3_2;
wire[15:0]    reg_weight21_4_1;
wire[15:0]    reg_psum21_4_1;
wire[15:0]    reg_weight21_4_2;
wire[15:0]    reg_psum21_4_2;
wire[15:0]    reg_weight21_5_1;
wire[15:0]    reg_psum21_5_1;
wire[15:0]    reg_weight21_5_2;
wire[15:0]    reg_psum21_5_2;
wire[15:0]    reg_weight21_6_1;
wire[15:0]    reg_psum21_6_1;
wire[15:0]    reg_weight21_6_2;
wire[15:0]    reg_psum21_6_2;
wire[15:0]    reg_weight21_7_1;
wire[15:0]    reg_psum21_7_1;
wire[15:0]    reg_weight21_7_2;
wire[15:0]    reg_psum21_7_2;
wire[15:0]    reg_weight21_8_1;
wire[15:0]    reg_psum21_8_1;
wire[15:0]    reg_weight21_8_2;
wire[15:0]    reg_psum21_8_2;
wire[15:0]    reg_weight21_9_1;
wire[15:0]    reg_psum21_9_1;
wire[15:0]    reg_weight21_9_2;
wire[15:0]    reg_psum21_9_2;
wire[15:0]    reg_weight21_10_1;
wire[15:0]    reg_psum21_10_1;
wire[15:0]    reg_weight21_10_2;
wire[15:0]    reg_psum21_10_2;
wire[15:0]    reg_weight21_11_1;
wire[15:0]    reg_psum21_11_1;
wire[15:0]    reg_weight21_11_2;
wire[15:0]    reg_psum21_11_2;
wire[15:0]    reg_weight21_12_1;
wire[15:0]    reg_psum21_12_1;
wire[15:0]    reg_weight21_12_2;
wire[15:0]    reg_psum21_12_2;
wire[15:0]    reg_weight21_13_1;
wire[15:0]    reg_psum21_13_1;
wire[15:0]    reg_weight21_13_2;
wire[15:0]    reg_psum21_13_2;
wire[15:0]    reg_weight21_14_1;
wire[15:0]    reg_psum21_14_1;
wire[15:0]    reg_weight21_14_2;
wire[15:0]    reg_psum21_14_2;
wire[15:0]    reg_weight21_15_1;
wire[15:0]    reg_psum21_15_1;
wire[15:0]    reg_weight21_15_2;
wire[15:0]    reg_psum21_15_2;
wire[15:0]    reg_weight21_16_1;
wire[15:0]    reg_psum21_16_1;
wire[15:0]    reg_weight21_16_2;
wire[15:0]    reg_psum21_16_2;
wire[15:0]    reg_weight21_17_1;
wire[15:0]    reg_psum21_17_1;
wire[15:0]    reg_weight21_17_2;
wire[15:0]    reg_psum21_17_2;
wire[15:0]    reg_weight21_18_1;
wire[15:0]    reg_psum21_18_1;
wire[15:0]    reg_weight21_18_2;
wire[15:0]    reg_psum21_18_2;
wire[15:0]    reg_weight21_19_1;
wire[15:0]    reg_psum21_19_1;
wire[15:0]    reg_weight21_19_2;
wire[15:0]    reg_psum21_19_2;
wire[15:0]    reg_weight21_20_1;
wire[15:0]    reg_psum21_20_1;
wire[15:0]    reg_weight21_20_2;
wire[15:0]    reg_psum21_20_2;
wire[15:0]    reg_weight21_21_1;
wire[15:0]    reg_psum21_21_1;
wire[15:0]    reg_weight21_21_2;
wire[15:0]    reg_psum21_21_2;
wire[15:0]    reg_weight21_22_1;
wire[15:0]    reg_psum21_22_1;
wire[15:0]    reg_weight21_22_2;
wire[15:0]    reg_psum21_22_2;
wire[15:0]    reg_weight21_23_1;
wire[15:0]    reg_psum21_23_1;
wire[15:0]    reg_weight21_23_2;
wire[15:0]    reg_psum21_23_2;
wire[15:0]    reg_weight21_24_1;
wire[15:0]    reg_psum21_24_1;
wire[15:0]    reg_weight21_24_2;
wire[15:0]    reg_psum21_24_2;
wire[15:0]    reg_weight21_25_1;
wire[15:0]    reg_psum21_25_1;
wire[15:0]    reg_weight21_25_2;
wire[15:0]    reg_psum21_25_2;
wire[15:0]    reg_weight21_26_1;
wire[15:0]    reg_psum21_26_1;
wire[15:0]    reg_weight21_26_2;
wire[15:0]    reg_psum21_26_2;
wire[15:0]    reg_weight21_27_1;
wire[15:0]    reg_psum21_27_1;
wire[15:0]    reg_weight21_27_2;
wire[15:0]    reg_psum21_27_2;
wire[15:0]    reg_weight21_28_1;
wire[15:0]    reg_psum21_28_1;
wire[15:0]    reg_weight21_28_2;
wire[15:0]    reg_psum21_28_2;
wire[15:0]    reg_weight21_29_1;
wire[15:0]    reg_psum21_29_1;
wire[15:0]    reg_weight21_29_2;
wire[15:0]    reg_psum21_29_2;
wire[15:0]    reg_weight21_30_1;
wire[15:0]    reg_psum21_30_1;
wire[15:0]    reg_weight21_30_2;
wire[15:0]    reg_psum21_30_2;
wire[15:0]    reg_weight21_31_1;
wire[15:0]    reg_psum21_31_1;
wire[15:0]    reg_weight21_31_2;
wire[15:0]    reg_psum21_31_2;
wire[15:0]    reg_weight21_32_1;
wire[15:0]    reg_psum21_32_1;
wire[15:0]    reg_weight21_32_2;
wire[15:0]    reg_psum21_32_2;
wire[15:0]    reg_weight22_1_1;
wire[15:0]    reg_psum22_1_1;
wire[15:0]    reg_weight22_1_2;
wire[15:0]    reg_psum22_1_2;
wire[15:0]    reg_weight22_2_1;
wire[15:0]    reg_psum22_2_1;
wire[15:0]    reg_weight22_2_2;
wire[15:0]    reg_psum22_2_2;
wire[15:0]    reg_weight22_3_1;
wire[15:0]    reg_psum22_3_1;
wire[15:0]    reg_weight22_3_2;
wire[15:0]    reg_psum22_3_2;
wire[15:0]    reg_weight22_4_1;
wire[15:0]    reg_psum22_4_1;
wire[15:0]    reg_weight22_4_2;
wire[15:0]    reg_psum22_4_2;
wire[15:0]    reg_weight22_5_1;
wire[15:0]    reg_psum22_5_1;
wire[15:0]    reg_weight22_5_2;
wire[15:0]    reg_psum22_5_2;
wire[15:0]    reg_weight22_6_1;
wire[15:0]    reg_psum22_6_1;
wire[15:0]    reg_weight22_6_2;
wire[15:0]    reg_psum22_6_2;
wire[15:0]    reg_weight22_7_1;
wire[15:0]    reg_psum22_7_1;
wire[15:0]    reg_weight22_7_2;
wire[15:0]    reg_psum22_7_2;
wire[15:0]    reg_weight22_8_1;
wire[15:0]    reg_psum22_8_1;
wire[15:0]    reg_weight22_8_2;
wire[15:0]    reg_psum22_8_2;
wire[15:0]    reg_weight22_9_1;
wire[15:0]    reg_psum22_9_1;
wire[15:0]    reg_weight22_9_2;
wire[15:0]    reg_psum22_9_2;
wire[15:0]    reg_weight22_10_1;
wire[15:0]    reg_psum22_10_1;
wire[15:0]    reg_weight22_10_2;
wire[15:0]    reg_psum22_10_2;
wire[15:0]    reg_weight22_11_1;
wire[15:0]    reg_psum22_11_1;
wire[15:0]    reg_weight22_11_2;
wire[15:0]    reg_psum22_11_2;
wire[15:0]    reg_weight22_12_1;
wire[15:0]    reg_psum22_12_1;
wire[15:0]    reg_weight22_12_2;
wire[15:0]    reg_psum22_12_2;
wire[15:0]    reg_weight22_13_1;
wire[15:0]    reg_psum22_13_1;
wire[15:0]    reg_weight22_13_2;
wire[15:0]    reg_psum22_13_2;
wire[15:0]    reg_weight22_14_1;
wire[15:0]    reg_psum22_14_1;
wire[15:0]    reg_weight22_14_2;
wire[15:0]    reg_psum22_14_2;
wire[15:0]    reg_weight22_15_1;
wire[15:0]    reg_psum22_15_1;
wire[15:0]    reg_weight22_15_2;
wire[15:0]    reg_psum22_15_2;
wire[15:0]    reg_weight22_16_1;
wire[15:0]    reg_psum22_16_1;
wire[15:0]    reg_weight22_16_2;
wire[15:0]    reg_psum22_16_2;
wire[15:0]    reg_weight22_17_1;
wire[15:0]    reg_psum22_17_1;
wire[15:0]    reg_weight22_17_2;
wire[15:0]    reg_psum22_17_2;
wire[15:0]    reg_weight22_18_1;
wire[15:0]    reg_psum22_18_1;
wire[15:0]    reg_weight22_18_2;
wire[15:0]    reg_psum22_18_2;
wire[15:0]    reg_weight22_19_1;
wire[15:0]    reg_psum22_19_1;
wire[15:0]    reg_weight22_19_2;
wire[15:0]    reg_psum22_19_2;
wire[15:0]    reg_weight22_20_1;
wire[15:0]    reg_psum22_20_1;
wire[15:0]    reg_weight22_20_2;
wire[15:0]    reg_psum22_20_2;
wire[15:0]    reg_weight22_21_1;
wire[15:0]    reg_psum22_21_1;
wire[15:0]    reg_weight22_21_2;
wire[15:0]    reg_psum22_21_2;
wire[15:0]    reg_weight22_22_1;
wire[15:0]    reg_psum22_22_1;
wire[15:0]    reg_weight22_22_2;
wire[15:0]    reg_psum22_22_2;
wire[15:0]    reg_weight22_23_1;
wire[15:0]    reg_psum22_23_1;
wire[15:0]    reg_weight22_23_2;
wire[15:0]    reg_psum22_23_2;
wire[15:0]    reg_weight22_24_1;
wire[15:0]    reg_psum22_24_1;
wire[15:0]    reg_weight22_24_2;
wire[15:0]    reg_psum22_24_2;
wire[15:0]    reg_weight22_25_1;
wire[15:0]    reg_psum22_25_1;
wire[15:0]    reg_weight22_25_2;
wire[15:0]    reg_psum22_25_2;
wire[15:0]    reg_weight22_26_1;
wire[15:0]    reg_psum22_26_1;
wire[15:0]    reg_weight22_26_2;
wire[15:0]    reg_psum22_26_2;
wire[15:0]    reg_weight22_27_1;
wire[15:0]    reg_psum22_27_1;
wire[15:0]    reg_weight22_27_2;
wire[15:0]    reg_psum22_27_2;
wire[15:0]    reg_weight22_28_1;
wire[15:0]    reg_psum22_28_1;
wire[15:0]    reg_weight22_28_2;
wire[15:0]    reg_psum22_28_2;
wire[15:0]    reg_weight22_29_1;
wire[15:0]    reg_psum22_29_1;
wire[15:0]    reg_weight22_29_2;
wire[15:0]    reg_psum22_29_2;
wire[15:0]    reg_weight22_30_1;
wire[15:0]    reg_psum22_30_1;
wire[15:0]    reg_weight22_30_2;
wire[15:0]    reg_psum22_30_2;
wire[15:0]    reg_weight22_31_1;
wire[15:0]    reg_psum22_31_1;
wire[15:0]    reg_weight22_31_2;
wire[15:0]    reg_psum22_31_2;
wire[15:0]    reg_weight22_32_1;
wire[15:0]    reg_psum22_32_1;
wire[15:0]    reg_weight22_32_2;
wire[15:0]    reg_psum22_32_2;
wire[15:0]    reg_weight23_1_1;
wire[15:0]    reg_psum23_1_1;
wire[15:0]    reg_weight23_1_2;
wire[15:0]    reg_psum23_1_2;
wire[15:0]    reg_weight23_2_1;
wire[15:0]    reg_psum23_2_1;
wire[15:0]    reg_weight23_2_2;
wire[15:0]    reg_psum23_2_2;
wire[15:0]    reg_weight23_3_1;
wire[15:0]    reg_psum23_3_1;
wire[15:0]    reg_weight23_3_2;
wire[15:0]    reg_psum23_3_2;
wire[15:0]    reg_weight23_4_1;
wire[15:0]    reg_psum23_4_1;
wire[15:0]    reg_weight23_4_2;
wire[15:0]    reg_psum23_4_2;
wire[15:0]    reg_weight23_5_1;
wire[15:0]    reg_psum23_5_1;
wire[15:0]    reg_weight23_5_2;
wire[15:0]    reg_psum23_5_2;
wire[15:0]    reg_weight23_6_1;
wire[15:0]    reg_psum23_6_1;
wire[15:0]    reg_weight23_6_2;
wire[15:0]    reg_psum23_6_2;
wire[15:0]    reg_weight23_7_1;
wire[15:0]    reg_psum23_7_1;
wire[15:0]    reg_weight23_7_2;
wire[15:0]    reg_psum23_7_2;
wire[15:0]    reg_weight23_8_1;
wire[15:0]    reg_psum23_8_1;
wire[15:0]    reg_weight23_8_2;
wire[15:0]    reg_psum23_8_2;
wire[15:0]    reg_weight23_9_1;
wire[15:0]    reg_psum23_9_1;
wire[15:0]    reg_weight23_9_2;
wire[15:0]    reg_psum23_9_2;
wire[15:0]    reg_weight23_10_1;
wire[15:0]    reg_psum23_10_1;
wire[15:0]    reg_weight23_10_2;
wire[15:0]    reg_psum23_10_2;
wire[15:0]    reg_weight23_11_1;
wire[15:0]    reg_psum23_11_1;
wire[15:0]    reg_weight23_11_2;
wire[15:0]    reg_psum23_11_2;
wire[15:0]    reg_weight23_12_1;
wire[15:0]    reg_psum23_12_1;
wire[15:0]    reg_weight23_12_2;
wire[15:0]    reg_psum23_12_2;
wire[15:0]    reg_weight23_13_1;
wire[15:0]    reg_psum23_13_1;
wire[15:0]    reg_weight23_13_2;
wire[15:0]    reg_psum23_13_2;
wire[15:0]    reg_weight23_14_1;
wire[15:0]    reg_psum23_14_1;
wire[15:0]    reg_weight23_14_2;
wire[15:0]    reg_psum23_14_2;
wire[15:0]    reg_weight23_15_1;
wire[15:0]    reg_psum23_15_1;
wire[15:0]    reg_weight23_15_2;
wire[15:0]    reg_psum23_15_2;
wire[15:0]    reg_weight23_16_1;
wire[15:0]    reg_psum23_16_1;
wire[15:0]    reg_weight23_16_2;
wire[15:0]    reg_psum23_16_2;
wire[15:0]    reg_weight23_17_1;
wire[15:0]    reg_psum23_17_1;
wire[15:0]    reg_weight23_17_2;
wire[15:0]    reg_psum23_17_2;
wire[15:0]    reg_weight23_18_1;
wire[15:0]    reg_psum23_18_1;
wire[15:0]    reg_weight23_18_2;
wire[15:0]    reg_psum23_18_2;
wire[15:0]    reg_weight23_19_1;
wire[15:0]    reg_psum23_19_1;
wire[15:0]    reg_weight23_19_2;
wire[15:0]    reg_psum23_19_2;
wire[15:0]    reg_weight23_20_1;
wire[15:0]    reg_psum23_20_1;
wire[15:0]    reg_weight23_20_2;
wire[15:0]    reg_psum23_20_2;
wire[15:0]    reg_weight23_21_1;
wire[15:0]    reg_psum23_21_1;
wire[15:0]    reg_weight23_21_2;
wire[15:0]    reg_psum23_21_2;
wire[15:0]    reg_weight23_22_1;
wire[15:0]    reg_psum23_22_1;
wire[15:0]    reg_weight23_22_2;
wire[15:0]    reg_psum23_22_2;
wire[15:0]    reg_weight23_23_1;
wire[15:0]    reg_psum23_23_1;
wire[15:0]    reg_weight23_23_2;
wire[15:0]    reg_psum23_23_2;
wire[15:0]    reg_weight23_24_1;
wire[15:0]    reg_psum23_24_1;
wire[15:0]    reg_weight23_24_2;
wire[15:0]    reg_psum23_24_2;
wire[15:0]    reg_weight23_25_1;
wire[15:0]    reg_psum23_25_1;
wire[15:0]    reg_weight23_25_2;
wire[15:0]    reg_psum23_25_2;
wire[15:0]    reg_weight23_26_1;
wire[15:0]    reg_psum23_26_1;
wire[15:0]    reg_weight23_26_2;
wire[15:0]    reg_psum23_26_2;
wire[15:0]    reg_weight23_27_1;
wire[15:0]    reg_psum23_27_1;
wire[15:0]    reg_weight23_27_2;
wire[15:0]    reg_psum23_27_2;
wire[15:0]    reg_weight23_28_1;
wire[15:0]    reg_psum23_28_1;
wire[15:0]    reg_weight23_28_2;
wire[15:0]    reg_psum23_28_2;
wire[15:0]    reg_weight23_29_1;
wire[15:0]    reg_psum23_29_1;
wire[15:0]    reg_weight23_29_2;
wire[15:0]    reg_psum23_29_2;
wire[15:0]    reg_weight23_30_1;
wire[15:0]    reg_psum23_30_1;
wire[15:0]    reg_weight23_30_2;
wire[15:0]    reg_psum23_30_2;
wire[15:0]    reg_weight23_31_1;
wire[15:0]    reg_psum23_31_1;
wire[15:0]    reg_weight23_31_2;
wire[15:0]    reg_psum23_31_2;
wire[15:0]    reg_weight23_32_1;
wire[15:0]    reg_psum23_32_1;
wire[15:0]    reg_weight23_32_2;
wire[15:0]    reg_psum23_32_2;
wire[15:0]    reg_weight24_1_1;
wire[15:0]    reg_psum24_1_1;
wire[15:0]    reg_weight24_1_2;
wire[15:0]    reg_psum24_1_2;
wire[15:0]    reg_weight24_2_1;
wire[15:0]    reg_psum24_2_1;
wire[15:0]    reg_weight24_2_2;
wire[15:0]    reg_psum24_2_2;
wire[15:0]    reg_weight24_3_1;
wire[15:0]    reg_psum24_3_1;
wire[15:0]    reg_weight24_3_2;
wire[15:0]    reg_psum24_3_2;
wire[15:0]    reg_weight24_4_1;
wire[15:0]    reg_psum24_4_1;
wire[15:0]    reg_weight24_4_2;
wire[15:0]    reg_psum24_4_2;
wire[15:0]    reg_weight24_5_1;
wire[15:0]    reg_psum24_5_1;
wire[15:0]    reg_weight24_5_2;
wire[15:0]    reg_psum24_5_2;
wire[15:0]    reg_weight24_6_1;
wire[15:0]    reg_psum24_6_1;
wire[15:0]    reg_weight24_6_2;
wire[15:0]    reg_psum24_6_2;
wire[15:0]    reg_weight24_7_1;
wire[15:0]    reg_psum24_7_1;
wire[15:0]    reg_weight24_7_2;
wire[15:0]    reg_psum24_7_2;
wire[15:0]    reg_weight24_8_1;
wire[15:0]    reg_psum24_8_1;
wire[15:0]    reg_weight24_8_2;
wire[15:0]    reg_psum24_8_2;
wire[15:0]    reg_weight24_9_1;
wire[15:0]    reg_psum24_9_1;
wire[15:0]    reg_weight24_9_2;
wire[15:0]    reg_psum24_9_2;
wire[15:0]    reg_weight24_10_1;
wire[15:0]    reg_psum24_10_1;
wire[15:0]    reg_weight24_10_2;
wire[15:0]    reg_psum24_10_2;
wire[15:0]    reg_weight24_11_1;
wire[15:0]    reg_psum24_11_1;
wire[15:0]    reg_weight24_11_2;
wire[15:0]    reg_psum24_11_2;
wire[15:0]    reg_weight24_12_1;
wire[15:0]    reg_psum24_12_1;
wire[15:0]    reg_weight24_12_2;
wire[15:0]    reg_psum24_12_2;
wire[15:0]    reg_weight24_13_1;
wire[15:0]    reg_psum24_13_1;
wire[15:0]    reg_weight24_13_2;
wire[15:0]    reg_psum24_13_2;
wire[15:0]    reg_weight24_14_1;
wire[15:0]    reg_psum24_14_1;
wire[15:0]    reg_weight24_14_2;
wire[15:0]    reg_psum24_14_2;
wire[15:0]    reg_weight24_15_1;
wire[15:0]    reg_psum24_15_1;
wire[15:0]    reg_weight24_15_2;
wire[15:0]    reg_psum24_15_2;
wire[15:0]    reg_weight24_16_1;
wire[15:0]    reg_psum24_16_1;
wire[15:0]    reg_weight24_16_2;
wire[15:0]    reg_psum24_16_2;
wire[15:0]    reg_weight24_17_1;
wire[15:0]    reg_psum24_17_1;
wire[15:0]    reg_weight24_17_2;
wire[15:0]    reg_psum24_17_2;
wire[15:0]    reg_weight24_18_1;
wire[15:0]    reg_psum24_18_1;
wire[15:0]    reg_weight24_18_2;
wire[15:0]    reg_psum24_18_2;
wire[15:0]    reg_weight24_19_1;
wire[15:0]    reg_psum24_19_1;
wire[15:0]    reg_weight24_19_2;
wire[15:0]    reg_psum24_19_2;
wire[15:0]    reg_weight24_20_1;
wire[15:0]    reg_psum24_20_1;
wire[15:0]    reg_weight24_20_2;
wire[15:0]    reg_psum24_20_2;
wire[15:0]    reg_weight24_21_1;
wire[15:0]    reg_psum24_21_1;
wire[15:0]    reg_weight24_21_2;
wire[15:0]    reg_psum24_21_2;
wire[15:0]    reg_weight24_22_1;
wire[15:0]    reg_psum24_22_1;
wire[15:0]    reg_weight24_22_2;
wire[15:0]    reg_psum24_22_2;
wire[15:0]    reg_weight24_23_1;
wire[15:0]    reg_psum24_23_1;
wire[15:0]    reg_weight24_23_2;
wire[15:0]    reg_psum24_23_2;
wire[15:0]    reg_weight24_24_1;
wire[15:0]    reg_psum24_24_1;
wire[15:0]    reg_weight24_24_2;
wire[15:0]    reg_psum24_24_2;
wire[15:0]    reg_weight24_25_1;
wire[15:0]    reg_psum24_25_1;
wire[15:0]    reg_weight24_25_2;
wire[15:0]    reg_psum24_25_2;
wire[15:0]    reg_weight24_26_1;
wire[15:0]    reg_psum24_26_1;
wire[15:0]    reg_weight24_26_2;
wire[15:0]    reg_psum24_26_2;
wire[15:0]    reg_weight24_27_1;
wire[15:0]    reg_psum24_27_1;
wire[15:0]    reg_weight24_27_2;
wire[15:0]    reg_psum24_27_2;
wire[15:0]    reg_weight24_28_1;
wire[15:0]    reg_psum24_28_1;
wire[15:0]    reg_weight24_28_2;
wire[15:0]    reg_psum24_28_2;
wire[15:0]    reg_weight24_29_1;
wire[15:0]    reg_psum24_29_1;
wire[15:0]    reg_weight24_29_2;
wire[15:0]    reg_psum24_29_2;
wire[15:0]    reg_weight24_30_1;
wire[15:0]    reg_psum24_30_1;
wire[15:0]    reg_weight24_30_2;
wire[15:0]    reg_psum24_30_2;
wire[15:0]    reg_weight24_31_1;
wire[15:0]    reg_psum24_31_1;
wire[15:0]    reg_weight24_31_2;
wire[15:0]    reg_psum24_31_2;
wire[15:0]    reg_weight24_32_1;
wire[15:0]    reg_psum24_32_1;
wire[15:0]    reg_weight24_32_2;
wire[15:0]    reg_psum24_32_2;
wire[15:0]    reg_weight25_1_1;
wire[15:0]    reg_psum25_1_1;
wire[15:0]    reg_weight25_1_2;
wire[15:0]    reg_psum25_1_2;
wire[15:0]    reg_weight25_2_1;
wire[15:0]    reg_psum25_2_1;
wire[15:0]    reg_weight25_2_2;
wire[15:0]    reg_psum25_2_2;
wire[15:0]    reg_weight25_3_1;
wire[15:0]    reg_psum25_3_1;
wire[15:0]    reg_weight25_3_2;
wire[15:0]    reg_psum25_3_2;
wire[15:0]    reg_weight25_4_1;
wire[15:0]    reg_psum25_4_1;
wire[15:0]    reg_weight25_4_2;
wire[15:0]    reg_psum25_4_2;
wire[15:0]    reg_weight25_5_1;
wire[15:0]    reg_psum25_5_1;
wire[15:0]    reg_weight25_5_2;
wire[15:0]    reg_psum25_5_2;
wire[15:0]    reg_weight25_6_1;
wire[15:0]    reg_psum25_6_1;
wire[15:0]    reg_weight25_6_2;
wire[15:0]    reg_psum25_6_2;
wire[15:0]    reg_weight25_7_1;
wire[15:0]    reg_psum25_7_1;
wire[15:0]    reg_weight25_7_2;
wire[15:0]    reg_psum25_7_2;
wire[15:0]    reg_weight25_8_1;
wire[15:0]    reg_psum25_8_1;
wire[15:0]    reg_weight25_8_2;
wire[15:0]    reg_psum25_8_2;
wire[15:0]    reg_weight25_9_1;
wire[15:0]    reg_psum25_9_1;
wire[15:0]    reg_weight25_9_2;
wire[15:0]    reg_psum25_9_2;
wire[15:0]    reg_weight25_10_1;
wire[15:0]    reg_psum25_10_1;
wire[15:0]    reg_weight25_10_2;
wire[15:0]    reg_psum25_10_2;
wire[15:0]    reg_weight25_11_1;
wire[15:0]    reg_psum25_11_1;
wire[15:0]    reg_weight25_11_2;
wire[15:0]    reg_psum25_11_2;
wire[15:0]    reg_weight25_12_1;
wire[15:0]    reg_psum25_12_1;
wire[15:0]    reg_weight25_12_2;
wire[15:0]    reg_psum25_12_2;
wire[15:0]    reg_weight25_13_1;
wire[15:0]    reg_psum25_13_1;
wire[15:0]    reg_weight25_13_2;
wire[15:0]    reg_psum25_13_2;
wire[15:0]    reg_weight25_14_1;
wire[15:0]    reg_psum25_14_1;
wire[15:0]    reg_weight25_14_2;
wire[15:0]    reg_psum25_14_2;
wire[15:0]    reg_weight25_15_1;
wire[15:0]    reg_psum25_15_1;
wire[15:0]    reg_weight25_15_2;
wire[15:0]    reg_psum25_15_2;
wire[15:0]    reg_weight25_16_1;
wire[15:0]    reg_psum25_16_1;
wire[15:0]    reg_weight25_16_2;
wire[15:0]    reg_psum25_16_2;
wire[15:0]    reg_weight25_17_1;
wire[15:0]    reg_psum25_17_1;
wire[15:0]    reg_weight25_17_2;
wire[15:0]    reg_psum25_17_2;
wire[15:0]    reg_weight25_18_1;
wire[15:0]    reg_psum25_18_1;
wire[15:0]    reg_weight25_18_2;
wire[15:0]    reg_psum25_18_2;
wire[15:0]    reg_weight25_19_1;
wire[15:0]    reg_psum25_19_1;
wire[15:0]    reg_weight25_19_2;
wire[15:0]    reg_psum25_19_2;
wire[15:0]    reg_weight25_20_1;
wire[15:0]    reg_psum25_20_1;
wire[15:0]    reg_weight25_20_2;
wire[15:0]    reg_psum25_20_2;
wire[15:0]    reg_weight25_21_1;
wire[15:0]    reg_psum25_21_1;
wire[15:0]    reg_weight25_21_2;
wire[15:0]    reg_psum25_21_2;
wire[15:0]    reg_weight25_22_1;
wire[15:0]    reg_psum25_22_1;
wire[15:0]    reg_weight25_22_2;
wire[15:0]    reg_psum25_22_2;
wire[15:0]    reg_weight25_23_1;
wire[15:0]    reg_psum25_23_1;
wire[15:0]    reg_weight25_23_2;
wire[15:0]    reg_psum25_23_2;
wire[15:0]    reg_weight25_24_1;
wire[15:0]    reg_psum25_24_1;
wire[15:0]    reg_weight25_24_2;
wire[15:0]    reg_psum25_24_2;
wire[15:0]    reg_weight25_25_1;
wire[15:0]    reg_psum25_25_1;
wire[15:0]    reg_weight25_25_2;
wire[15:0]    reg_psum25_25_2;
wire[15:0]    reg_weight25_26_1;
wire[15:0]    reg_psum25_26_1;
wire[15:0]    reg_weight25_26_2;
wire[15:0]    reg_psum25_26_2;
wire[15:0]    reg_weight25_27_1;
wire[15:0]    reg_psum25_27_1;
wire[15:0]    reg_weight25_27_2;
wire[15:0]    reg_psum25_27_2;
wire[15:0]    reg_weight25_28_1;
wire[15:0]    reg_psum25_28_1;
wire[15:0]    reg_weight25_28_2;
wire[15:0]    reg_psum25_28_2;
wire[15:0]    reg_weight25_29_1;
wire[15:0]    reg_psum25_29_1;
wire[15:0]    reg_weight25_29_2;
wire[15:0]    reg_psum25_29_2;
wire[15:0]    reg_weight25_30_1;
wire[15:0]    reg_psum25_30_1;
wire[15:0]    reg_weight25_30_2;
wire[15:0]    reg_psum25_30_2;
wire[15:0]    reg_weight25_31_1;
wire[15:0]    reg_psum25_31_1;
wire[15:0]    reg_weight25_31_2;
wire[15:0]    reg_psum25_31_2;
wire[15:0]    reg_weight25_32_1;
wire[15:0]    reg_psum25_32_1;
wire[15:0]    reg_weight25_32_2;
wire[15:0]    reg_psum25_32_2;
wire[15:0]    reg_weight26_1_1;
wire[15:0]    reg_psum26_1_1;
wire[15:0]    reg_weight26_1_2;
wire[15:0]    reg_psum26_1_2;
wire[15:0]    reg_weight26_2_1;
wire[15:0]    reg_psum26_2_1;
wire[15:0]    reg_weight26_2_2;
wire[15:0]    reg_psum26_2_2;
wire[15:0]    reg_weight26_3_1;
wire[15:0]    reg_psum26_3_1;
wire[15:0]    reg_weight26_3_2;
wire[15:0]    reg_psum26_3_2;
wire[15:0]    reg_weight26_4_1;
wire[15:0]    reg_psum26_4_1;
wire[15:0]    reg_weight26_4_2;
wire[15:0]    reg_psum26_4_2;
wire[15:0]    reg_weight26_5_1;
wire[15:0]    reg_psum26_5_1;
wire[15:0]    reg_weight26_5_2;
wire[15:0]    reg_psum26_5_2;
wire[15:0]    reg_weight26_6_1;
wire[15:0]    reg_psum26_6_1;
wire[15:0]    reg_weight26_6_2;
wire[15:0]    reg_psum26_6_2;
wire[15:0]    reg_weight26_7_1;
wire[15:0]    reg_psum26_7_1;
wire[15:0]    reg_weight26_7_2;
wire[15:0]    reg_psum26_7_2;
wire[15:0]    reg_weight26_8_1;
wire[15:0]    reg_psum26_8_1;
wire[15:0]    reg_weight26_8_2;
wire[15:0]    reg_psum26_8_2;
wire[15:0]    reg_weight26_9_1;
wire[15:0]    reg_psum26_9_1;
wire[15:0]    reg_weight26_9_2;
wire[15:0]    reg_psum26_9_2;
wire[15:0]    reg_weight26_10_1;
wire[15:0]    reg_psum26_10_1;
wire[15:0]    reg_weight26_10_2;
wire[15:0]    reg_psum26_10_2;
wire[15:0]    reg_weight26_11_1;
wire[15:0]    reg_psum26_11_1;
wire[15:0]    reg_weight26_11_2;
wire[15:0]    reg_psum26_11_2;
wire[15:0]    reg_weight26_12_1;
wire[15:0]    reg_psum26_12_1;
wire[15:0]    reg_weight26_12_2;
wire[15:0]    reg_psum26_12_2;
wire[15:0]    reg_weight26_13_1;
wire[15:0]    reg_psum26_13_1;
wire[15:0]    reg_weight26_13_2;
wire[15:0]    reg_psum26_13_2;
wire[15:0]    reg_weight26_14_1;
wire[15:0]    reg_psum26_14_1;
wire[15:0]    reg_weight26_14_2;
wire[15:0]    reg_psum26_14_2;
wire[15:0]    reg_weight26_15_1;
wire[15:0]    reg_psum26_15_1;
wire[15:0]    reg_weight26_15_2;
wire[15:0]    reg_psum26_15_2;
wire[15:0]    reg_weight26_16_1;
wire[15:0]    reg_psum26_16_1;
wire[15:0]    reg_weight26_16_2;
wire[15:0]    reg_psum26_16_2;
wire[15:0]    reg_weight26_17_1;
wire[15:0]    reg_psum26_17_1;
wire[15:0]    reg_weight26_17_2;
wire[15:0]    reg_psum26_17_2;
wire[15:0]    reg_weight26_18_1;
wire[15:0]    reg_psum26_18_1;
wire[15:0]    reg_weight26_18_2;
wire[15:0]    reg_psum26_18_2;
wire[15:0]    reg_weight26_19_1;
wire[15:0]    reg_psum26_19_1;
wire[15:0]    reg_weight26_19_2;
wire[15:0]    reg_psum26_19_2;
wire[15:0]    reg_weight26_20_1;
wire[15:0]    reg_psum26_20_1;
wire[15:0]    reg_weight26_20_2;
wire[15:0]    reg_psum26_20_2;
wire[15:0]    reg_weight26_21_1;
wire[15:0]    reg_psum26_21_1;
wire[15:0]    reg_weight26_21_2;
wire[15:0]    reg_psum26_21_2;
wire[15:0]    reg_weight26_22_1;
wire[15:0]    reg_psum26_22_1;
wire[15:0]    reg_weight26_22_2;
wire[15:0]    reg_psum26_22_2;
wire[15:0]    reg_weight26_23_1;
wire[15:0]    reg_psum26_23_1;
wire[15:0]    reg_weight26_23_2;
wire[15:0]    reg_psum26_23_2;
wire[15:0]    reg_weight26_24_1;
wire[15:0]    reg_psum26_24_1;
wire[15:0]    reg_weight26_24_2;
wire[15:0]    reg_psum26_24_2;
wire[15:0]    reg_weight26_25_1;
wire[15:0]    reg_psum26_25_1;
wire[15:0]    reg_weight26_25_2;
wire[15:0]    reg_psum26_25_2;
wire[15:0]    reg_weight26_26_1;
wire[15:0]    reg_psum26_26_1;
wire[15:0]    reg_weight26_26_2;
wire[15:0]    reg_psum26_26_2;
wire[15:0]    reg_weight26_27_1;
wire[15:0]    reg_psum26_27_1;
wire[15:0]    reg_weight26_27_2;
wire[15:0]    reg_psum26_27_2;
wire[15:0]    reg_weight26_28_1;
wire[15:0]    reg_psum26_28_1;
wire[15:0]    reg_weight26_28_2;
wire[15:0]    reg_psum26_28_2;
wire[15:0]    reg_weight26_29_1;
wire[15:0]    reg_psum26_29_1;
wire[15:0]    reg_weight26_29_2;
wire[15:0]    reg_psum26_29_2;
wire[15:0]    reg_weight26_30_1;
wire[15:0]    reg_psum26_30_1;
wire[15:0]    reg_weight26_30_2;
wire[15:0]    reg_psum26_30_2;
wire[15:0]    reg_weight26_31_1;
wire[15:0]    reg_psum26_31_1;
wire[15:0]    reg_weight26_31_2;
wire[15:0]    reg_psum26_31_2;
wire[15:0]    reg_weight26_32_1;
wire[15:0]    reg_psum26_32_1;
wire[15:0]    reg_weight26_32_2;
wire[15:0]    reg_psum26_32_2;
wire[15:0]    reg_weight27_1_1;
wire[15:0]    reg_psum27_1_1;
wire[15:0]    reg_weight27_1_2;
wire[15:0]    reg_psum27_1_2;
wire[15:0]    reg_weight27_2_1;
wire[15:0]    reg_psum27_2_1;
wire[15:0]    reg_weight27_2_2;
wire[15:0]    reg_psum27_2_2;
wire[15:0]    reg_weight27_3_1;
wire[15:0]    reg_psum27_3_1;
wire[15:0]    reg_weight27_3_2;
wire[15:0]    reg_psum27_3_2;
wire[15:0]    reg_weight27_4_1;
wire[15:0]    reg_psum27_4_1;
wire[15:0]    reg_weight27_4_2;
wire[15:0]    reg_psum27_4_2;
wire[15:0]    reg_weight27_5_1;
wire[15:0]    reg_psum27_5_1;
wire[15:0]    reg_weight27_5_2;
wire[15:0]    reg_psum27_5_2;
wire[15:0]    reg_weight27_6_1;
wire[15:0]    reg_psum27_6_1;
wire[15:0]    reg_weight27_6_2;
wire[15:0]    reg_psum27_6_2;
wire[15:0]    reg_weight27_7_1;
wire[15:0]    reg_psum27_7_1;
wire[15:0]    reg_weight27_7_2;
wire[15:0]    reg_psum27_7_2;
wire[15:0]    reg_weight27_8_1;
wire[15:0]    reg_psum27_8_1;
wire[15:0]    reg_weight27_8_2;
wire[15:0]    reg_psum27_8_2;
wire[15:0]    reg_weight27_9_1;
wire[15:0]    reg_psum27_9_1;
wire[15:0]    reg_weight27_9_2;
wire[15:0]    reg_psum27_9_2;
wire[15:0]    reg_weight27_10_1;
wire[15:0]    reg_psum27_10_1;
wire[15:0]    reg_weight27_10_2;
wire[15:0]    reg_psum27_10_2;
wire[15:0]    reg_weight27_11_1;
wire[15:0]    reg_psum27_11_1;
wire[15:0]    reg_weight27_11_2;
wire[15:0]    reg_psum27_11_2;
wire[15:0]    reg_weight27_12_1;
wire[15:0]    reg_psum27_12_1;
wire[15:0]    reg_weight27_12_2;
wire[15:0]    reg_psum27_12_2;
wire[15:0]    reg_weight27_13_1;
wire[15:0]    reg_psum27_13_1;
wire[15:0]    reg_weight27_13_2;
wire[15:0]    reg_psum27_13_2;
wire[15:0]    reg_weight27_14_1;
wire[15:0]    reg_psum27_14_1;
wire[15:0]    reg_weight27_14_2;
wire[15:0]    reg_psum27_14_2;
wire[15:0]    reg_weight27_15_1;
wire[15:0]    reg_psum27_15_1;
wire[15:0]    reg_weight27_15_2;
wire[15:0]    reg_psum27_15_2;
wire[15:0]    reg_weight27_16_1;
wire[15:0]    reg_psum27_16_1;
wire[15:0]    reg_weight27_16_2;
wire[15:0]    reg_psum27_16_2;
wire[15:0]    reg_weight27_17_1;
wire[15:0]    reg_psum27_17_1;
wire[15:0]    reg_weight27_17_2;
wire[15:0]    reg_psum27_17_2;
wire[15:0]    reg_weight27_18_1;
wire[15:0]    reg_psum27_18_1;
wire[15:0]    reg_weight27_18_2;
wire[15:0]    reg_psum27_18_2;
wire[15:0]    reg_weight27_19_1;
wire[15:0]    reg_psum27_19_1;
wire[15:0]    reg_weight27_19_2;
wire[15:0]    reg_psum27_19_2;
wire[15:0]    reg_weight27_20_1;
wire[15:0]    reg_psum27_20_1;
wire[15:0]    reg_weight27_20_2;
wire[15:0]    reg_psum27_20_2;
wire[15:0]    reg_weight27_21_1;
wire[15:0]    reg_psum27_21_1;
wire[15:0]    reg_weight27_21_2;
wire[15:0]    reg_psum27_21_2;
wire[15:0]    reg_weight27_22_1;
wire[15:0]    reg_psum27_22_1;
wire[15:0]    reg_weight27_22_2;
wire[15:0]    reg_psum27_22_2;
wire[15:0]    reg_weight27_23_1;
wire[15:0]    reg_psum27_23_1;
wire[15:0]    reg_weight27_23_2;
wire[15:0]    reg_psum27_23_2;
wire[15:0]    reg_weight27_24_1;
wire[15:0]    reg_psum27_24_1;
wire[15:0]    reg_weight27_24_2;
wire[15:0]    reg_psum27_24_2;
wire[15:0]    reg_weight27_25_1;
wire[15:0]    reg_psum27_25_1;
wire[15:0]    reg_weight27_25_2;
wire[15:0]    reg_psum27_25_2;
wire[15:0]    reg_weight27_26_1;
wire[15:0]    reg_psum27_26_1;
wire[15:0]    reg_weight27_26_2;
wire[15:0]    reg_psum27_26_2;
wire[15:0]    reg_weight27_27_1;
wire[15:0]    reg_psum27_27_1;
wire[15:0]    reg_weight27_27_2;
wire[15:0]    reg_psum27_27_2;
wire[15:0]    reg_weight27_28_1;
wire[15:0]    reg_psum27_28_1;
wire[15:0]    reg_weight27_28_2;
wire[15:0]    reg_psum27_28_2;
wire[15:0]    reg_weight27_29_1;
wire[15:0]    reg_psum27_29_1;
wire[15:0]    reg_weight27_29_2;
wire[15:0]    reg_psum27_29_2;
wire[15:0]    reg_weight27_30_1;
wire[15:0]    reg_psum27_30_1;
wire[15:0]    reg_weight27_30_2;
wire[15:0]    reg_psum27_30_2;
wire[15:0]    reg_weight27_31_1;
wire[15:0]    reg_psum27_31_1;
wire[15:0]    reg_weight27_31_2;
wire[15:0]    reg_psum27_31_2;
wire[15:0]    reg_weight27_32_1;
wire[15:0]    reg_psum27_32_1;
wire[15:0]    reg_weight27_32_2;
wire[15:0]    reg_psum27_32_2;
wire[15:0]    reg_weight28_1_1;
wire[15:0]    reg_psum28_1_1;
wire[15:0]    reg_weight28_1_2;
wire[15:0]    reg_psum28_1_2;
wire[15:0]    reg_weight28_2_1;
wire[15:0]    reg_psum28_2_1;
wire[15:0]    reg_weight28_2_2;
wire[15:0]    reg_psum28_2_2;
wire[15:0]    reg_weight28_3_1;
wire[15:0]    reg_psum28_3_1;
wire[15:0]    reg_weight28_3_2;
wire[15:0]    reg_psum28_3_2;
wire[15:0]    reg_weight28_4_1;
wire[15:0]    reg_psum28_4_1;
wire[15:0]    reg_weight28_4_2;
wire[15:0]    reg_psum28_4_2;
wire[15:0]    reg_weight28_5_1;
wire[15:0]    reg_psum28_5_1;
wire[15:0]    reg_weight28_5_2;
wire[15:0]    reg_psum28_5_2;
wire[15:0]    reg_weight28_6_1;
wire[15:0]    reg_psum28_6_1;
wire[15:0]    reg_weight28_6_2;
wire[15:0]    reg_psum28_6_2;
wire[15:0]    reg_weight28_7_1;
wire[15:0]    reg_psum28_7_1;
wire[15:0]    reg_weight28_7_2;
wire[15:0]    reg_psum28_7_2;
wire[15:0]    reg_weight28_8_1;
wire[15:0]    reg_psum28_8_1;
wire[15:0]    reg_weight28_8_2;
wire[15:0]    reg_psum28_8_2;
wire[15:0]    reg_weight28_9_1;
wire[15:0]    reg_psum28_9_1;
wire[15:0]    reg_weight28_9_2;
wire[15:0]    reg_psum28_9_2;
wire[15:0]    reg_weight28_10_1;
wire[15:0]    reg_psum28_10_1;
wire[15:0]    reg_weight28_10_2;
wire[15:0]    reg_psum28_10_2;
wire[15:0]    reg_weight28_11_1;
wire[15:0]    reg_psum28_11_1;
wire[15:0]    reg_weight28_11_2;
wire[15:0]    reg_psum28_11_2;
wire[15:0]    reg_weight28_12_1;
wire[15:0]    reg_psum28_12_1;
wire[15:0]    reg_weight28_12_2;
wire[15:0]    reg_psum28_12_2;
wire[15:0]    reg_weight28_13_1;
wire[15:0]    reg_psum28_13_1;
wire[15:0]    reg_weight28_13_2;
wire[15:0]    reg_psum28_13_2;
wire[15:0]    reg_weight28_14_1;
wire[15:0]    reg_psum28_14_1;
wire[15:0]    reg_weight28_14_2;
wire[15:0]    reg_psum28_14_2;
wire[15:0]    reg_weight28_15_1;
wire[15:0]    reg_psum28_15_1;
wire[15:0]    reg_weight28_15_2;
wire[15:0]    reg_psum28_15_2;
wire[15:0]    reg_weight28_16_1;
wire[15:0]    reg_psum28_16_1;
wire[15:0]    reg_weight28_16_2;
wire[15:0]    reg_psum28_16_2;
wire[15:0]    reg_weight28_17_1;
wire[15:0]    reg_psum28_17_1;
wire[15:0]    reg_weight28_17_2;
wire[15:0]    reg_psum28_17_2;
wire[15:0]    reg_weight28_18_1;
wire[15:0]    reg_psum28_18_1;
wire[15:0]    reg_weight28_18_2;
wire[15:0]    reg_psum28_18_2;
wire[15:0]    reg_weight28_19_1;
wire[15:0]    reg_psum28_19_1;
wire[15:0]    reg_weight28_19_2;
wire[15:0]    reg_psum28_19_2;
wire[15:0]    reg_weight28_20_1;
wire[15:0]    reg_psum28_20_1;
wire[15:0]    reg_weight28_20_2;
wire[15:0]    reg_psum28_20_2;
wire[15:0]    reg_weight28_21_1;
wire[15:0]    reg_psum28_21_1;
wire[15:0]    reg_weight28_21_2;
wire[15:0]    reg_psum28_21_2;
wire[15:0]    reg_weight28_22_1;
wire[15:0]    reg_psum28_22_1;
wire[15:0]    reg_weight28_22_2;
wire[15:0]    reg_psum28_22_2;
wire[15:0]    reg_weight28_23_1;
wire[15:0]    reg_psum28_23_1;
wire[15:0]    reg_weight28_23_2;
wire[15:0]    reg_psum28_23_2;
wire[15:0]    reg_weight28_24_1;
wire[15:0]    reg_psum28_24_1;
wire[15:0]    reg_weight28_24_2;
wire[15:0]    reg_psum28_24_2;
wire[15:0]    reg_weight28_25_1;
wire[15:0]    reg_psum28_25_1;
wire[15:0]    reg_weight28_25_2;
wire[15:0]    reg_psum28_25_2;
wire[15:0]    reg_weight28_26_1;
wire[15:0]    reg_psum28_26_1;
wire[15:0]    reg_weight28_26_2;
wire[15:0]    reg_psum28_26_2;
wire[15:0]    reg_weight28_27_1;
wire[15:0]    reg_psum28_27_1;
wire[15:0]    reg_weight28_27_2;
wire[15:0]    reg_psum28_27_2;
wire[15:0]    reg_weight28_28_1;
wire[15:0]    reg_psum28_28_1;
wire[15:0]    reg_weight28_28_2;
wire[15:0]    reg_psum28_28_2;
wire[15:0]    reg_weight28_29_1;
wire[15:0]    reg_psum28_29_1;
wire[15:0]    reg_weight28_29_2;
wire[15:0]    reg_psum28_29_2;
wire[15:0]    reg_weight28_30_1;
wire[15:0]    reg_psum28_30_1;
wire[15:0]    reg_weight28_30_2;
wire[15:0]    reg_psum28_30_2;
wire[15:0]    reg_weight28_31_1;
wire[15:0]    reg_psum28_31_1;
wire[15:0]    reg_weight28_31_2;
wire[15:0]    reg_psum28_31_2;
wire[15:0]    reg_weight28_32_1;
wire[15:0]    reg_psum28_32_1;
wire[15:0]    reg_weight28_32_2;
wire[15:0]    reg_psum28_32_2;
wire[15:0]    reg_weight29_1_1;
wire[15:0]    reg_psum29_1_1;
wire[15:0]    reg_weight29_1_2;
wire[15:0]    reg_psum29_1_2;
wire[15:0]    reg_weight29_2_1;
wire[15:0]    reg_psum29_2_1;
wire[15:0]    reg_weight29_2_2;
wire[15:0]    reg_psum29_2_2;
wire[15:0]    reg_weight29_3_1;
wire[15:0]    reg_psum29_3_1;
wire[15:0]    reg_weight29_3_2;
wire[15:0]    reg_psum29_3_2;
wire[15:0]    reg_weight29_4_1;
wire[15:0]    reg_psum29_4_1;
wire[15:0]    reg_weight29_4_2;
wire[15:0]    reg_psum29_4_2;
wire[15:0]    reg_weight29_5_1;
wire[15:0]    reg_psum29_5_1;
wire[15:0]    reg_weight29_5_2;
wire[15:0]    reg_psum29_5_2;
wire[15:0]    reg_weight29_6_1;
wire[15:0]    reg_psum29_6_1;
wire[15:0]    reg_weight29_6_2;
wire[15:0]    reg_psum29_6_2;
wire[15:0]    reg_weight29_7_1;
wire[15:0]    reg_psum29_7_1;
wire[15:0]    reg_weight29_7_2;
wire[15:0]    reg_psum29_7_2;
wire[15:0]    reg_weight29_8_1;
wire[15:0]    reg_psum29_8_1;
wire[15:0]    reg_weight29_8_2;
wire[15:0]    reg_psum29_8_2;
wire[15:0]    reg_weight29_9_1;
wire[15:0]    reg_psum29_9_1;
wire[15:0]    reg_weight29_9_2;
wire[15:0]    reg_psum29_9_2;
wire[15:0]    reg_weight29_10_1;
wire[15:0]    reg_psum29_10_1;
wire[15:0]    reg_weight29_10_2;
wire[15:0]    reg_psum29_10_2;
wire[15:0]    reg_weight29_11_1;
wire[15:0]    reg_psum29_11_1;
wire[15:0]    reg_weight29_11_2;
wire[15:0]    reg_psum29_11_2;
wire[15:0]    reg_weight29_12_1;
wire[15:0]    reg_psum29_12_1;
wire[15:0]    reg_weight29_12_2;
wire[15:0]    reg_psum29_12_2;
wire[15:0]    reg_weight29_13_1;
wire[15:0]    reg_psum29_13_1;
wire[15:0]    reg_weight29_13_2;
wire[15:0]    reg_psum29_13_2;
wire[15:0]    reg_weight29_14_1;
wire[15:0]    reg_psum29_14_1;
wire[15:0]    reg_weight29_14_2;
wire[15:0]    reg_psum29_14_2;
wire[15:0]    reg_weight29_15_1;
wire[15:0]    reg_psum29_15_1;
wire[15:0]    reg_weight29_15_2;
wire[15:0]    reg_psum29_15_2;
wire[15:0]    reg_weight29_16_1;
wire[15:0]    reg_psum29_16_1;
wire[15:0]    reg_weight29_16_2;
wire[15:0]    reg_psum29_16_2;
wire[15:0]    reg_weight29_17_1;
wire[15:0]    reg_psum29_17_1;
wire[15:0]    reg_weight29_17_2;
wire[15:0]    reg_psum29_17_2;
wire[15:0]    reg_weight29_18_1;
wire[15:0]    reg_psum29_18_1;
wire[15:0]    reg_weight29_18_2;
wire[15:0]    reg_psum29_18_2;
wire[15:0]    reg_weight29_19_1;
wire[15:0]    reg_psum29_19_1;
wire[15:0]    reg_weight29_19_2;
wire[15:0]    reg_psum29_19_2;
wire[15:0]    reg_weight29_20_1;
wire[15:0]    reg_psum29_20_1;
wire[15:0]    reg_weight29_20_2;
wire[15:0]    reg_psum29_20_2;
wire[15:0]    reg_weight29_21_1;
wire[15:0]    reg_psum29_21_1;
wire[15:0]    reg_weight29_21_2;
wire[15:0]    reg_psum29_21_2;
wire[15:0]    reg_weight29_22_1;
wire[15:0]    reg_psum29_22_1;
wire[15:0]    reg_weight29_22_2;
wire[15:0]    reg_psum29_22_2;
wire[15:0]    reg_weight29_23_1;
wire[15:0]    reg_psum29_23_1;
wire[15:0]    reg_weight29_23_2;
wire[15:0]    reg_psum29_23_2;
wire[15:0]    reg_weight29_24_1;
wire[15:0]    reg_psum29_24_1;
wire[15:0]    reg_weight29_24_2;
wire[15:0]    reg_psum29_24_2;
wire[15:0]    reg_weight29_25_1;
wire[15:0]    reg_psum29_25_1;
wire[15:0]    reg_weight29_25_2;
wire[15:0]    reg_psum29_25_2;
wire[15:0]    reg_weight29_26_1;
wire[15:0]    reg_psum29_26_1;
wire[15:0]    reg_weight29_26_2;
wire[15:0]    reg_psum29_26_2;
wire[15:0]    reg_weight29_27_1;
wire[15:0]    reg_psum29_27_1;
wire[15:0]    reg_weight29_27_2;
wire[15:0]    reg_psum29_27_2;
wire[15:0]    reg_weight29_28_1;
wire[15:0]    reg_psum29_28_1;
wire[15:0]    reg_weight29_28_2;
wire[15:0]    reg_psum29_28_2;
wire[15:0]    reg_weight29_29_1;
wire[15:0]    reg_psum29_29_1;
wire[15:0]    reg_weight29_29_2;
wire[15:0]    reg_psum29_29_2;
wire[15:0]    reg_weight29_30_1;
wire[15:0]    reg_psum29_30_1;
wire[15:0]    reg_weight29_30_2;
wire[15:0]    reg_psum29_30_2;
wire[15:0]    reg_weight29_31_1;
wire[15:0]    reg_psum29_31_1;
wire[15:0]    reg_weight29_31_2;
wire[15:0]    reg_psum29_31_2;
wire[15:0]    reg_weight29_32_1;
wire[15:0]    reg_psum29_32_1;
wire[15:0]    reg_weight29_32_2;
wire[15:0]    reg_psum29_32_2;
wire[15:0]    reg_weight30_1_1;
wire[15:0]    reg_psum30_1_1;
wire[15:0]    reg_weight30_1_2;
wire[15:0]    reg_psum30_1_2;
wire[15:0]    reg_weight30_2_1;
wire[15:0]    reg_psum30_2_1;
wire[15:0]    reg_weight30_2_2;
wire[15:0]    reg_psum30_2_2;
wire[15:0]    reg_weight30_3_1;
wire[15:0]    reg_psum30_3_1;
wire[15:0]    reg_weight30_3_2;
wire[15:0]    reg_psum30_3_2;
wire[15:0]    reg_weight30_4_1;
wire[15:0]    reg_psum30_4_1;
wire[15:0]    reg_weight30_4_2;
wire[15:0]    reg_psum30_4_2;
wire[15:0]    reg_weight30_5_1;
wire[15:0]    reg_psum30_5_1;
wire[15:0]    reg_weight30_5_2;
wire[15:0]    reg_psum30_5_2;
wire[15:0]    reg_weight30_6_1;
wire[15:0]    reg_psum30_6_1;
wire[15:0]    reg_weight30_6_2;
wire[15:0]    reg_psum30_6_2;
wire[15:0]    reg_weight30_7_1;
wire[15:0]    reg_psum30_7_1;
wire[15:0]    reg_weight30_7_2;
wire[15:0]    reg_psum30_7_2;
wire[15:0]    reg_weight30_8_1;
wire[15:0]    reg_psum30_8_1;
wire[15:0]    reg_weight30_8_2;
wire[15:0]    reg_psum30_8_2;
wire[15:0]    reg_weight30_9_1;
wire[15:0]    reg_psum30_9_1;
wire[15:0]    reg_weight30_9_2;
wire[15:0]    reg_psum30_9_2;
wire[15:0]    reg_weight30_10_1;
wire[15:0]    reg_psum30_10_1;
wire[15:0]    reg_weight30_10_2;
wire[15:0]    reg_psum30_10_2;
wire[15:0]    reg_weight30_11_1;
wire[15:0]    reg_psum30_11_1;
wire[15:0]    reg_weight30_11_2;
wire[15:0]    reg_psum30_11_2;
wire[15:0]    reg_weight30_12_1;
wire[15:0]    reg_psum30_12_1;
wire[15:0]    reg_weight30_12_2;
wire[15:0]    reg_psum30_12_2;
wire[15:0]    reg_weight30_13_1;
wire[15:0]    reg_psum30_13_1;
wire[15:0]    reg_weight30_13_2;
wire[15:0]    reg_psum30_13_2;
wire[15:0]    reg_weight30_14_1;
wire[15:0]    reg_psum30_14_1;
wire[15:0]    reg_weight30_14_2;
wire[15:0]    reg_psum30_14_2;
wire[15:0]    reg_weight30_15_1;
wire[15:0]    reg_psum30_15_1;
wire[15:0]    reg_weight30_15_2;
wire[15:0]    reg_psum30_15_2;
wire[15:0]    reg_weight30_16_1;
wire[15:0]    reg_psum30_16_1;
wire[15:0]    reg_weight30_16_2;
wire[15:0]    reg_psum30_16_2;
wire[15:0]    reg_weight30_17_1;
wire[15:0]    reg_psum30_17_1;
wire[15:0]    reg_weight30_17_2;
wire[15:0]    reg_psum30_17_2;
wire[15:0]    reg_weight30_18_1;
wire[15:0]    reg_psum30_18_1;
wire[15:0]    reg_weight30_18_2;
wire[15:0]    reg_psum30_18_2;
wire[15:0]    reg_weight30_19_1;
wire[15:0]    reg_psum30_19_1;
wire[15:0]    reg_weight30_19_2;
wire[15:0]    reg_psum30_19_2;
wire[15:0]    reg_weight30_20_1;
wire[15:0]    reg_psum30_20_1;
wire[15:0]    reg_weight30_20_2;
wire[15:0]    reg_psum30_20_2;
wire[15:0]    reg_weight30_21_1;
wire[15:0]    reg_psum30_21_1;
wire[15:0]    reg_weight30_21_2;
wire[15:0]    reg_psum30_21_2;
wire[15:0]    reg_weight30_22_1;
wire[15:0]    reg_psum30_22_1;
wire[15:0]    reg_weight30_22_2;
wire[15:0]    reg_psum30_22_2;
wire[15:0]    reg_weight30_23_1;
wire[15:0]    reg_psum30_23_1;
wire[15:0]    reg_weight30_23_2;
wire[15:0]    reg_psum30_23_2;
wire[15:0]    reg_weight30_24_1;
wire[15:0]    reg_psum30_24_1;
wire[15:0]    reg_weight30_24_2;
wire[15:0]    reg_psum30_24_2;
wire[15:0]    reg_weight30_25_1;
wire[15:0]    reg_psum30_25_1;
wire[15:0]    reg_weight30_25_2;
wire[15:0]    reg_psum30_25_2;
wire[15:0]    reg_weight30_26_1;
wire[15:0]    reg_psum30_26_1;
wire[15:0]    reg_weight30_26_2;
wire[15:0]    reg_psum30_26_2;
wire[15:0]    reg_weight30_27_1;
wire[15:0]    reg_psum30_27_1;
wire[15:0]    reg_weight30_27_2;
wire[15:0]    reg_psum30_27_2;
wire[15:0]    reg_weight30_28_1;
wire[15:0]    reg_psum30_28_1;
wire[15:0]    reg_weight30_28_2;
wire[15:0]    reg_psum30_28_2;
wire[15:0]    reg_weight30_29_1;
wire[15:0]    reg_psum30_29_1;
wire[15:0]    reg_weight30_29_2;
wire[15:0]    reg_psum30_29_2;
wire[15:0]    reg_weight30_30_1;
wire[15:0]    reg_psum30_30_1;
wire[15:0]    reg_weight30_30_2;
wire[15:0]    reg_psum30_30_2;
wire[15:0]    reg_weight30_31_1;
wire[15:0]    reg_psum30_31_1;
wire[15:0]    reg_weight30_31_2;
wire[15:0]    reg_psum30_31_2;
wire[15:0]    reg_weight30_32_1;
wire[15:0]    reg_psum30_32_1;
wire[15:0]    reg_weight30_32_2;
wire[15:0]    reg_psum30_32_2;
wire[15:0]    reg_weight31_1_1;
wire[15:0]    reg_psum31_1_1;
wire[15:0]    reg_weight31_1_2;
wire[15:0]    reg_psum31_1_2;
wire[15:0]    reg_weight31_2_1;
wire[15:0]    reg_psum31_2_1;
wire[15:0]    reg_weight31_2_2;
wire[15:0]    reg_psum31_2_2;
wire[15:0]    reg_weight31_3_1;
wire[15:0]    reg_psum31_3_1;
wire[15:0]    reg_weight31_3_2;
wire[15:0]    reg_psum31_3_2;
wire[15:0]    reg_weight31_4_1;
wire[15:0]    reg_psum31_4_1;
wire[15:0]    reg_weight31_4_2;
wire[15:0]    reg_psum31_4_2;
wire[15:0]    reg_weight31_5_1;
wire[15:0]    reg_psum31_5_1;
wire[15:0]    reg_weight31_5_2;
wire[15:0]    reg_psum31_5_2;
wire[15:0]    reg_weight31_6_1;
wire[15:0]    reg_psum31_6_1;
wire[15:0]    reg_weight31_6_2;
wire[15:0]    reg_psum31_6_2;
wire[15:0]    reg_weight31_7_1;
wire[15:0]    reg_psum31_7_1;
wire[15:0]    reg_weight31_7_2;
wire[15:0]    reg_psum31_7_2;
wire[15:0]    reg_weight31_8_1;
wire[15:0]    reg_psum31_8_1;
wire[15:0]    reg_weight31_8_2;
wire[15:0]    reg_psum31_8_2;
wire[15:0]    reg_weight31_9_1;
wire[15:0]    reg_psum31_9_1;
wire[15:0]    reg_weight31_9_2;
wire[15:0]    reg_psum31_9_2;
wire[15:0]    reg_weight31_10_1;
wire[15:0]    reg_psum31_10_1;
wire[15:0]    reg_weight31_10_2;
wire[15:0]    reg_psum31_10_2;
wire[15:0]    reg_weight31_11_1;
wire[15:0]    reg_psum31_11_1;
wire[15:0]    reg_weight31_11_2;
wire[15:0]    reg_psum31_11_2;
wire[15:0]    reg_weight31_12_1;
wire[15:0]    reg_psum31_12_1;
wire[15:0]    reg_weight31_12_2;
wire[15:0]    reg_psum31_12_2;
wire[15:0]    reg_weight31_13_1;
wire[15:0]    reg_psum31_13_1;
wire[15:0]    reg_weight31_13_2;
wire[15:0]    reg_psum31_13_2;
wire[15:0]    reg_weight31_14_1;
wire[15:0]    reg_psum31_14_1;
wire[15:0]    reg_weight31_14_2;
wire[15:0]    reg_psum31_14_2;
wire[15:0]    reg_weight31_15_1;
wire[15:0]    reg_psum31_15_1;
wire[15:0]    reg_weight31_15_2;
wire[15:0]    reg_psum31_15_2;
wire[15:0]    reg_weight31_16_1;
wire[15:0]    reg_psum31_16_1;
wire[15:0]    reg_weight31_16_2;
wire[15:0]    reg_psum31_16_2;
wire[15:0]    reg_weight31_17_1;
wire[15:0]    reg_psum31_17_1;
wire[15:0]    reg_weight31_17_2;
wire[15:0]    reg_psum31_17_2;
wire[15:0]    reg_weight31_18_1;
wire[15:0]    reg_psum31_18_1;
wire[15:0]    reg_weight31_18_2;
wire[15:0]    reg_psum31_18_2;
wire[15:0]    reg_weight31_19_1;
wire[15:0]    reg_psum31_19_1;
wire[15:0]    reg_weight31_19_2;
wire[15:0]    reg_psum31_19_2;
wire[15:0]    reg_weight31_20_1;
wire[15:0]    reg_psum31_20_1;
wire[15:0]    reg_weight31_20_2;
wire[15:0]    reg_psum31_20_2;
wire[15:0]    reg_weight31_21_1;
wire[15:0]    reg_psum31_21_1;
wire[15:0]    reg_weight31_21_2;
wire[15:0]    reg_psum31_21_2;
wire[15:0]    reg_weight31_22_1;
wire[15:0]    reg_psum31_22_1;
wire[15:0]    reg_weight31_22_2;
wire[15:0]    reg_psum31_22_2;
wire[15:0]    reg_weight31_23_1;
wire[15:0]    reg_psum31_23_1;
wire[15:0]    reg_weight31_23_2;
wire[15:0]    reg_psum31_23_2;
wire[15:0]    reg_weight31_24_1;
wire[15:0]    reg_psum31_24_1;
wire[15:0]    reg_weight31_24_2;
wire[15:0]    reg_psum31_24_2;
wire[15:0]    reg_weight31_25_1;
wire[15:0]    reg_psum31_25_1;
wire[15:0]    reg_weight31_25_2;
wire[15:0]    reg_psum31_25_2;
wire[15:0]    reg_weight31_26_1;
wire[15:0]    reg_psum31_26_1;
wire[15:0]    reg_weight31_26_2;
wire[15:0]    reg_psum31_26_2;
wire[15:0]    reg_weight31_27_1;
wire[15:0]    reg_psum31_27_1;
wire[15:0]    reg_weight31_27_2;
wire[15:0]    reg_psum31_27_2;
wire[15:0]    reg_weight31_28_1;
wire[15:0]    reg_psum31_28_1;
wire[15:0]    reg_weight31_28_2;
wire[15:0]    reg_psum31_28_2;
wire[15:0]    reg_weight31_29_1;
wire[15:0]    reg_psum31_29_1;
wire[15:0]    reg_weight31_29_2;
wire[15:0]    reg_psum31_29_2;
wire[15:0]    reg_weight31_30_1;
wire[15:0]    reg_psum31_30_1;
wire[15:0]    reg_weight31_30_2;
wire[15:0]    reg_psum31_30_2;
wire[15:0]    reg_weight31_31_1;
wire[15:0]    reg_psum31_31_1;
wire[15:0]    reg_weight31_31_2;
wire[15:0]    reg_psum31_31_2;
wire[15:0]    reg_weight31_32_1;
wire[15:0]    reg_psum31_32_1;
wire[15:0]    reg_weight31_32_2;
wire[15:0]    reg_psum31_32_2;
SA22 U1_1(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_1_1), .partial_sum_in12(in_psum1_1_2), .weight_in11(in_weight1_1_1), .weight_in12(in_weight1_1_2), .activation_in11(in_activation1_1_1), .activation_in21(in_activation1_1_2), .reg_partial_sum21(reg_psum1_1_1), .reg_partial_sum22(reg_psum1_1_2), .reg_weight21(reg_weight1_1_1), .reg_weight22(reg_weight1_1_2), .reg_activation12(reg_activation1_1_1), .reg_activation22(reg_activation1_1_2), .weight_en(weight_en));
SA22 U1_2(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_2_1), .partial_sum_in12(in_psum1_2_2), .weight_in11(in_weight1_2_1), .weight_in12(in_weight1_2_2), .activation_in11(reg_activation1_1_1), .activation_in21(reg_activation1_1_2), .reg_partial_sum21(reg_psum1_2_1), .reg_partial_sum22(reg_psum1_2_2), .reg_weight21(reg_weight1_2_1), .reg_weight22(reg_weight1_2_2), .reg_activation12(reg_activation1_2_1), .reg_activation22(reg_activation1_2_2), .weight_en(weight_en));
SA22 U1_3(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_3_1), .partial_sum_in12(in_psum1_3_2), .weight_in11(in_weight1_3_1), .weight_in12(in_weight1_3_2), .activation_in11(reg_activation1_2_1), .activation_in21(reg_activation1_2_2), .reg_partial_sum21(reg_psum1_3_1), .reg_partial_sum22(reg_psum1_3_2), .reg_weight21(reg_weight1_3_1), .reg_weight22(reg_weight1_3_2), .reg_activation12(reg_activation1_3_1), .reg_activation22(reg_activation1_3_2), .weight_en(weight_en));
SA22 U1_4(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_4_1), .partial_sum_in12(in_psum1_4_2), .weight_in11(in_weight1_4_1), .weight_in12(in_weight1_4_2), .activation_in11(reg_activation1_3_1), .activation_in21(reg_activation1_3_2), .reg_partial_sum21(reg_psum1_4_1), .reg_partial_sum22(reg_psum1_4_2), .reg_weight21(reg_weight1_4_1), .reg_weight22(reg_weight1_4_2), .reg_activation12(reg_activation1_4_1), .reg_activation22(reg_activation1_4_2), .weight_en(weight_en));
SA22 U1_5(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_5_1), .partial_sum_in12(in_psum1_5_2), .weight_in11(in_weight1_5_1), .weight_in12(in_weight1_5_2), .activation_in11(reg_activation1_4_1), .activation_in21(reg_activation1_4_2), .reg_partial_sum21(reg_psum1_5_1), .reg_partial_sum22(reg_psum1_5_2), .reg_weight21(reg_weight1_5_1), .reg_weight22(reg_weight1_5_2), .reg_activation12(reg_activation1_5_1), .reg_activation22(reg_activation1_5_2), .weight_en(weight_en));
SA22 U1_6(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_6_1), .partial_sum_in12(in_psum1_6_2), .weight_in11(in_weight1_6_1), .weight_in12(in_weight1_6_2), .activation_in11(reg_activation1_5_1), .activation_in21(reg_activation1_5_2), .reg_partial_sum21(reg_psum1_6_1), .reg_partial_sum22(reg_psum1_6_2), .reg_weight21(reg_weight1_6_1), .reg_weight22(reg_weight1_6_2), .reg_activation12(reg_activation1_6_1), .reg_activation22(reg_activation1_6_2), .weight_en(weight_en));
SA22 U1_7(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_7_1), .partial_sum_in12(in_psum1_7_2), .weight_in11(in_weight1_7_1), .weight_in12(in_weight1_7_2), .activation_in11(reg_activation1_6_1), .activation_in21(reg_activation1_6_2), .reg_partial_sum21(reg_psum1_7_1), .reg_partial_sum22(reg_psum1_7_2), .reg_weight21(reg_weight1_7_1), .reg_weight22(reg_weight1_7_2), .reg_activation12(reg_activation1_7_1), .reg_activation22(reg_activation1_7_2), .weight_en(weight_en));
SA22 U1_8(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_8_1), .partial_sum_in12(in_psum1_8_2), .weight_in11(in_weight1_8_1), .weight_in12(in_weight1_8_2), .activation_in11(reg_activation1_7_1), .activation_in21(reg_activation1_7_2), .reg_partial_sum21(reg_psum1_8_1), .reg_partial_sum22(reg_psum1_8_2), .reg_weight21(reg_weight1_8_1), .reg_weight22(reg_weight1_8_2), .reg_activation12(reg_activation1_8_1), .reg_activation22(reg_activation1_8_2), .weight_en(weight_en));
SA22 U1_9(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_9_1), .partial_sum_in12(in_psum1_9_2), .weight_in11(in_weight1_9_1), .weight_in12(in_weight1_9_2), .activation_in11(reg_activation1_8_1), .activation_in21(reg_activation1_8_2), .reg_partial_sum21(reg_psum1_9_1), .reg_partial_sum22(reg_psum1_9_2), .reg_weight21(reg_weight1_9_1), .reg_weight22(reg_weight1_9_2), .reg_activation12(reg_activation1_9_1), .reg_activation22(reg_activation1_9_2), .weight_en(weight_en));
SA22 U1_10(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_10_1), .partial_sum_in12(in_psum1_10_2), .weight_in11(in_weight1_10_1), .weight_in12(in_weight1_10_2), .activation_in11(reg_activation1_9_1), .activation_in21(reg_activation1_9_2), .reg_partial_sum21(reg_psum1_10_1), .reg_partial_sum22(reg_psum1_10_2), .reg_weight21(reg_weight1_10_1), .reg_weight22(reg_weight1_10_2), .reg_activation12(reg_activation1_10_1), .reg_activation22(reg_activation1_10_2), .weight_en(weight_en));
SA22 U1_11(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_11_1), .partial_sum_in12(in_psum1_11_2), .weight_in11(in_weight1_11_1), .weight_in12(in_weight1_11_2), .activation_in11(reg_activation1_10_1), .activation_in21(reg_activation1_10_2), .reg_partial_sum21(reg_psum1_11_1), .reg_partial_sum22(reg_psum1_11_2), .reg_weight21(reg_weight1_11_1), .reg_weight22(reg_weight1_11_2), .reg_activation12(reg_activation1_11_1), .reg_activation22(reg_activation1_11_2), .weight_en(weight_en));
SA22 U1_12(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_12_1), .partial_sum_in12(in_psum1_12_2), .weight_in11(in_weight1_12_1), .weight_in12(in_weight1_12_2), .activation_in11(reg_activation1_11_1), .activation_in21(reg_activation1_11_2), .reg_partial_sum21(reg_psum1_12_1), .reg_partial_sum22(reg_psum1_12_2), .reg_weight21(reg_weight1_12_1), .reg_weight22(reg_weight1_12_2), .reg_activation12(reg_activation1_12_1), .reg_activation22(reg_activation1_12_2), .weight_en(weight_en));
SA22 U1_13(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_13_1), .partial_sum_in12(in_psum1_13_2), .weight_in11(in_weight1_13_1), .weight_in12(in_weight1_13_2), .activation_in11(reg_activation1_12_1), .activation_in21(reg_activation1_12_2), .reg_partial_sum21(reg_psum1_13_1), .reg_partial_sum22(reg_psum1_13_2), .reg_weight21(reg_weight1_13_1), .reg_weight22(reg_weight1_13_2), .reg_activation12(reg_activation1_13_1), .reg_activation22(reg_activation1_13_2), .weight_en(weight_en));
SA22 U1_14(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_14_1), .partial_sum_in12(in_psum1_14_2), .weight_in11(in_weight1_14_1), .weight_in12(in_weight1_14_2), .activation_in11(reg_activation1_13_1), .activation_in21(reg_activation1_13_2), .reg_partial_sum21(reg_psum1_14_1), .reg_partial_sum22(reg_psum1_14_2), .reg_weight21(reg_weight1_14_1), .reg_weight22(reg_weight1_14_2), .reg_activation12(reg_activation1_14_1), .reg_activation22(reg_activation1_14_2), .weight_en(weight_en));
SA22 U1_15(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_15_1), .partial_sum_in12(in_psum1_15_2), .weight_in11(in_weight1_15_1), .weight_in12(in_weight1_15_2), .activation_in11(reg_activation1_14_1), .activation_in21(reg_activation1_14_2), .reg_partial_sum21(reg_psum1_15_1), .reg_partial_sum22(reg_psum1_15_2), .reg_weight21(reg_weight1_15_1), .reg_weight22(reg_weight1_15_2), .reg_activation12(reg_activation1_15_1), .reg_activation22(reg_activation1_15_2), .weight_en(weight_en));
SA22 U1_16(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_16_1), .partial_sum_in12(in_psum1_16_2), .weight_in11(in_weight1_16_1), .weight_in12(in_weight1_16_2), .activation_in11(reg_activation1_15_1), .activation_in21(reg_activation1_15_2), .reg_partial_sum21(reg_psum1_16_1), .reg_partial_sum22(reg_psum1_16_2), .reg_weight21(reg_weight1_16_1), .reg_weight22(reg_weight1_16_2), .reg_activation12(reg_activation1_16_1), .reg_activation22(reg_activation1_16_2), .weight_en(weight_en));
SA22 U1_17(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_17_1), .partial_sum_in12(in_psum1_17_2), .weight_in11(in_weight1_17_1), .weight_in12(in_weight1_17_2), .activation_in11(reg_activation1_16_1), .activation_in21(reg_activation1_16_2), .reg_partial_sum21(reg_psum1_17_1), .reg_partial_sum22(reg_psum1_17_2), .reg_weight21(reg_weight1_17_1), .reg_weight22(reg_weight1_17_2), .reg_activation12(reg_activation1_17_1), .reg_activation22(reg_activation1_17_2), .weight_en(weight_en));
SA22 U1_18(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_18_1), .partial_sum_in12(in_psum1_18_2), .weight_in11(in_weight1_18_1), .weight_in12(in_weight1_18_2), .activation_in11(reg_activation1_17_1), .activation_in21(reg_activation1_17_2), .reg_partial_sum21(reg_psum1_18_1), .reg_partial_sum22(reg_psum1_18_2), .reg_weight21(reg_weight1_18_1), .reg_weight22(reg_weight1_18_2), .reg_activation12(reg_activation1_18_1), .reg_activation22(reg_activation1_18_2), .weight_en(weight_en));
SA22 U1_19(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_19_1), .partial_sum_in12(in_psum1_19_2), .weight_in11(in_weight1_19_1), .weight_in12(in_weight1_19_2), .activation_in11(reg_activation1_18_1), .activation_in21(reg_activation1_18_2), .reg_partial_sum21(reg_psum1_19_1), .reg_partial_sum22(reg_psum1_19_2), .reg_weight21(reg_weight1_19_1), .reg_weight22(reg_weight1_19_2), .reg_activation12(reg_activation1_19_1), .reg_activation22(reg_activation1_19_2), .weight_en(weight_en));
SA22 U1_20(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_20_1), .partial_sum_in12(in_psum1_20_2), .weight_in11(in_weight1_20_1), .weight_in12(in_weight1_20_2), .activation_in11(reg_activation1_19_1), .activation_in21(reg_activation1_19_2), .reg_partial_sum21(reg_psum1_20_1), .reg_partial_sum22(reg_psum1_20_2), .reg_weight21(reg_weight1_20_1), .reg_weight22(reg_weight1_20_2), .reg_activation12(reg_activation1_20_1), .reg_activation22(reg_activation1_20_2), .weight_en(weight_en));
SA22 U1_21(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_21_1), .partial_sum_in12(in_psum1_21_2), .weight_in11(in_weight1_21_1), .weight_in12(in_weight1_21_2), .activation_in11(reg_activation1_20_1), .activation_in21(reg_activation1_20_2), .reg_partial_sum21(reg_psum1_21_1), .reg_partial_sum22(reg_psum1_21_2), .reg_weight21(reg_weight1_21_1), .reg_weight22(reg_weight1_21_2), .reg_activation12(reg_activation1_21_1), .reg_activation22(reg_activation1_21_2), .weight_en(weight_en));
SA22 U1_22(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_22_1), .partial_sum_in12(in_psum1_22_2), .weight_in11(in_weight1_22_1), .weight_in12(in_weight1_22_2), .activation_in11(reg_activation1_21_1), .activation_in21(reg_activation1_21_2), .reg_partial_sum21(reg_psum1_22_1), .reg_partial_sum22(reg_psum1_22_2), .reg_weight21(reg_weight1_22_1), .reg_weight22(reg_weight1_22_2), .reg_activation12(reg_activation1_22_1), .reg_activation22(reg_activation1_22_2), .weight_en(weight_en));
SA22 U1_23(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_23_1), .partial_sum_in12(in_psum1_23_2), .weight_in11(in_weight1_23_1), .weight_in12(in_weight1_23_2), .activation_in11(reg_activation1_22_1), .activation_in21(reg_activation1_22_2), .reg_partial_sum21(reg_psum1_23_1), .reg_partial_sum22(reg_psum1_23_2), .reg_weight21(reg_weight1_23_1), .reg_weight22(reg_weight1_23_2), .reg_activation12(reg_activation1_23_1), .reg_activation22(reg_activation1_23_2), .weight_en(weight_en));
SA22 U1_24(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_24_1), .partial_sum_in12(in_psum1_24_2), .weight_in11(in_weight1_24_1), .weight_in12(in_weight1_24_2), .activation_in11(reg_activation1_23_1), .activation_in21(reg_activation1_23_2), .reg_partial_sum21(reg_psum1_24_1), .reg_partial_sum22(reg_psum1_24_2), .reg_weight21(reg_weight1_24_1), .reg_weight22(reg_weight1_24_2), .reg_activation12(reg_activation1_24_1), .reg_activation22(reg_activation1_24_2), .weight_en(weight_en));
SA22 U1_25(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_25_1), .partial_sum_in12(in_psum1_25_2), .weight_in11(in_weight1_25_1), .weight_in12(in_weight1_25_2), .activation_in11(reg_activation1_24_1), .activation_in21(reg_activation1_24_2), .reg_partial_sum21(reg_psum1_25_1), .reg_partial_sum22(reg_psum1_25_2), .reg_weight21(reg_weight1_25_1), .reg_weight22(reg_weight1_25_2), .reg_activation12(reg_activation1_25_1), .reg_activation22(reg_activation1_25_2), .weight_en(weight_en));
SA22 U1_26(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_26_1), .partial_sum_in12(in_psum1_26_2), .weight_in11(in_weight1_26_1), .weight_in12(in_weight1_26_2), .activation_in11(reg_activation1_25_1), .activation_in21(reg_activation1_25_2), .reg_partial_sum21(reg_psum1_26_1), .reg_partial_sum22(reg_psum1_26_2), .reg_weight21(reg_weight1_26_1), .reg_weight22(reg_weight1_26_2), .reg_activation12(reg_activation1_26_1), .reg_activation22(reg_activation1_26_2), .weight_en(weight_en));
SA22 U1_27(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_27_1), .partial_sum_in12(in_psum1_27_2), .weight_in11(in_weight1_27_1), .weight_in12(in_weight1_27_2), .activation_in11(reg_activation1_26_1), .activation_in21(reg_activation1_26_2), .reg_partial_sum21(reg_psum1_27_1), .reg_partial_sum22(reg_psum1_27_2), .reg_weight21(reg_weight1_27_1), .reg_weight22(reg_weight1_27_2), .reg_activation12(reg_activation1_27_1), .reg_activation22(reg_activation1_27_2), .weight_en(weight_en));
SA22 U1_28(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_28_1), .partial_sum_in12(in_psum1_28_2), .weight_in11(in_weight1_28_1), .weight_in12(in_weight1_28_2), .activation_in11(reg_activation1_27_1), .activation_in21(reg_activation1_27_2), .reg_partial_sum21(reg_psum1_28_1), .reg_partial_sum22(reg_psum1_28_2), .reg_weight21(reg_weight1_28_1), .reg_weight22(reg_weight1_28_2), .reg_activation12(reg_activation1_28_1), .reg_activation22(reg_activation1_28_2), .weight_en(weight_en));
SA22 U1_29(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_29_1), .partial_sum_in12(in_psum1_29_2), .weight_in11(in_weight1_29_1), .weight_in12(in_weight1_29_2), .activation_in11(reg_activation1_28_1), .activation_in21(reg_activation1_28_2), .reg_partial_sum21(reg_psum1_29_1), .reg_partial_sum22(reg_psum1_29_2), .reg_weight21(reg_weight1_29_1), .reg_weight22(reg_weight1_29_2), .reg_activation12(reg_activation1_29_1), .reg_activation22(reg_activation1_29_2), .weight_en(weight_en));
SA22 U1_30(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_30_1), .partial_sum_in12(in_psum1_30_2), .weight_in11(in_weight1_30_1), .weight_in12(in_weight1_30_2), .activation_in11(reg_activation1_29_1), .activation_in21(reg_activation1_29_2), .reg_partial_sum21(reg_psum1_30_1), .reg_partial_sum22(reg_psum1_30_2), .reg_weight21(reg_weight1_30_1), .reg_weight22(reg_weight1_30_2), .reg_activation12(reg_activation1_30_1), .reg_activation22(reg_activation1_30_2), .weight_en(weight_en));
SA22 U1_31(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_31_1), .partial_sum_in12(in_psum1_31_2), .weight_in11(in_weight1_31_1), .weight_in12(in_weight1_31_2), .activation_in11(reg_activation1_30_1), .activation_in21(reg_activation1_30_2), .reg_partial_sum21(reg_psum1_31_1), .reg_partial_sum22(reg_psum1_31_2), .reg_weight21(reg_weight1_31_1), .reg_weight22(reg_weight1_31_2), .reg_activation12(reg_activation1_31_1), .reg_activation22(reg_activation1_31_2), .weight_en(weight_en));
SA22 U1_32(.clk(clk), .rst(rst), .partial_sum_in11(in_psum1_32_1), .partial_sum_in12(in_psum1_32_2), .weight_in11(in_weight1_32_1), .weight_in12(in_weight1_32_2), .activation_in11(reg_activation1_31_1), .activation_in21(reg_activation1_31_2), .reg_partial_sum21(reg_psum1_32_1), .reg_partial_sum22(reg_psum1_32_2), .reg_weight21(reg_weight1_32_1), .reg_weight22(reg_weight1_32_2), .weight_en(weight_en));
SA22 U2_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_1_1), .partial_sum_in12(reg_psum1_1_2), .weight_in11(reg_weight1_1_1), .weight_in12(reg_weight1_1_2), .activation_in11(in_activation2_1_1), .activation_in21(in_activation2_1_2), .reg_partial_sum21(reg_psum2_1_1), .reg_partial_sum22(reg_psum2_1_2), .reg_weight21(reg_weight2_1_1), .reg_weight22(reg_weight2_1_2), .reg_activation12(reg_activation2_1_1), .reg_activation22(reg_activation2_1_2), .weight_en(weight_en));
SA22 U2_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_2_1), .partial_sum_in12(reg_psum1_2_2), .weight_in11(reg_weight1_2_1), .weight_in12(reg_weight1_2_2), .activation_in11(reg_activation2_1_1), .activation_in21(reg_activation2_1_2), .reg_partial_sum21(reg_psum2_2_1), .reg_partial_sum22(reg_psum2_2_2), .reg_weight21(reg_weight2_2_1), .reg_weight22(reg_weight2_2_2), .reg_activation12(reg_activation2_2_1), .reg_activation22(reg_activation2_2_2), .weight_en(weight_en));
SA22 U2_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_3_1), .partial_sum_in12(reg_psum1_3_2), .weight_in11(reg_weight1_3_1), .weight_in12(reg_weight1_3_2), .activation_in11(reg_activation2_2_1), .activation_in21(reg_activation2_2_2), .reg_partial_sum21(reg_psum2_3_1), .reg_partial_sum22(reg_psum2_3_2), .reg_weight21(reg_weight2_3_1), .reg_weight22(reg_weight2_3_2), .reg_activation12(reg_activation2_3_1), .reg_activation22(reg_activation2_3_2), .weight_en(weight_en));
SA22 U2_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_4_1), .partial_sum_in12(reg_psum1_4_2), .weight_in11(reg_weight1_4_1), .weight_in12(reg_weight1_4_2), .activation_in11(reg_activation2_3_1), .activation_in21(reg_activation2_3_2), .reg_partial_sum21(reg_psum2_4_1), .reg_partial_sum22(reg_psum2_4_2), .reg_weight21(reg_weight2_4_1), .reg_weight22(reg_weight2_4_2), .reg_activation12(reg_activation2_4_1), .reg_activation22(reg_activation2_4_2), .weight_en(weight_en));
SA22 U2_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_5_1), .partial_sum_in12(reg_psum1_5_2), .weight_in11(reg_weight1_5_1), .weight_in12(reg_weight1_5_2), .activation_in11(reg_activation2_4_1), .activation_in21(reg_activation2_4_2), .reg_partial_sum21(reg_psum2_5_1), .reg_partial_sum22(reg_psum2_5_2), .reg_weight21(reg_weight2_5_1), .reg_weight22(reg_weight2_5_2), .reg_activation12(reg_activation2_5_1), .reg_activation22(reg_activation2_5_2), .weight_en(weight_en));
SA22 U2_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_6_1), .partial_sum_in12(reg_psum1_6_2), .weight_in11(reg_weight1_6_1), .weight_in12(reg_weight1_6_2), .activation_in11(reg_activation2_5_1), .activation_in21(reg_activation2_5_2), .reg_partial_sum21(reg_psum2_6_1), .reg_partial_sum22(reg_psum2_6_2), .reg_weight21(reg_weight2_6_1), .reg_weight22(reg_weight2_6_2), .reg_activation12(reg_activation2_6_1), .reg_activation22(reg_activation2_6_2), .weight_en(weight_en));
SA22 U2_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_7_1), .partial_sum_in12(reg_psum1_7_2), .weight_in11(reg_weight1_7_1), .weight_in12(reg_weight1_7_2), .activation_in11(reg_activation2_6_1), .activation_in21(reg_activation2_6_2), .reg_partial_sum21(reg_psum2_7_1), .reg_partial_sum22(reg_psum2_7_2), .reg_weight21(reg_weight2_7_1), .reg_weight22(reg_weight2_7_2), .reg_activation12(reg_activation2_7_1), .reg_activation22(reg_activation2_7_2), .weight_en(weight_en));
SA22 U2_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_8_1), .partial_sum_in12(reg_psum1_8_2), .weight_in11(reg_weight1_8_1), .weight_in12(reg_weight1_8_2), .activation_in11(reg_activation2_7_1), .activation_in21(reg_activation2_7_2), .reg_partial_sum21(reg_psum2_8_1), .reg_partial_sum22(reg_psum2_8_2), .reg_weight21(reg_weight2_8_1), .reg_weight22(reg_weight2_8_2), .reg_activation12(reg_activation2_8_1), .reg_activation22(reg_activation2_8_2), .weight_en(weight_en));
SA22 U2_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_9_1), .partial_sum_in12(reg_psum1_9_2), .weight_in11(reg_weight1_9_1), .weight_in12(reg_weight1_9_2), .activation_in11(reg_activation2_8_1), .activation_in21(reg_activation2_8_2), .reg_partial_sum21(reg_psum2_9_1), .reg_partial_sum22(reg_psum2_9_2), .reg_weight21(reg_weight2_9_1), .reg_weight22(reg_weight2_9_2), .reg_activation12(reg_activation2_9_1), .reg_activation22(reg_activation2_9_2), .weight_en(weight_en));
SA22 U2_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_10_1), .partial_sum_in12(reg_psum1_10_2), .weight_in11(reg_weight1_10_1), .weight_in12(reg_weight1_10_2), .activation_in11(reg_activation2_9_1), .activation_in21(reg_activation2_9_2), .reg_partial_sum21(reg_psum2_10_1), .reg_partial_sum22(reg_psum2_10_2), .reg_weight21(reg_weight2_10_1), .reg_weight22(reg_weight2_10_2), .reg_activation12(reg_activation2_10_1), .reg_activation22(reg_activation2_10_2), .weight_en(weight_en));
SA22 U2_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_11_1), .partial_sum_in12(reg_psum1_11_2), .weight_in11(reg_weight1_11_1), .weight_in12(reg_weight1_11_2), .activation_in11(reg_activation2_10_1), .activation_in21(reg_activation2_10_2), .reg_partial_sum21(reg_psum2_11_1), .reg_partial_sum22(reg_psum2_11_2), .reg_weight21(reg_weight2_11_1), .reg_weight22(reg_weight2_11_2), .reg_activation12(reg_activation2_11_1), .reg_activation22(reg_activation2_11_2), .weight_en(weight_en));
SA22 U2_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_12_1), .partial_sum_in12(reg_psum1_12_2), .weight_in11(reg_weight1_12_1), .weight_in12(reg_weight1_12_2), .activation_in11(reg_activation2_11_1), .activation_in21(reg_activation2_11_2), .reg_partial_sum21(reg_psum2_12_1), .reg_partial_sum22(reg_psum2_12_2), .reg_weight21(reg_weight2_12_1), .reg_weight22(reg_weight2_12_2), .reg_activation12(reg_activation2_12_1), .reg_activation22(reg_activation2_12_2), .weight_en(weight_en));
SA22 U2_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_13_1), .partial_sum_in12(reg_psum1_13_2), .weight_in11(reg_weight1_13_1), .weight_in12(reg_weight1_13_2), .activation_in11(reg_activation2_12_1), .activation_in21(reg_activation2_12_2), .reg_partial_sum21(reg_psum2_13_1), .reg_partial_sum22(reg_psum2_13_2), .reg_weight21(reg_weight2_13_1), .reg_weight22(reg_weight2_13_2), .reg_activation12(reg_activation2_13_1), .reg_activation22(reg_activation2_13_2), .weight_en(weight_en));
SA22 U2_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_14_1), .partial_sum_in12(reg_psum1_14_2), .weight_in11(reg_weight1_14_1), .weight_in12(reg_weight1_14_2), .activation_in11(reg_activation2_13_1), .activation_in21(reg_activation2_13_2), .reg_partial_sum21(reg_psum2_14_1), .reg_partial_sum22(reg_psum2_14_2), .reg_weight21(reg_weight2_14_1), .reg_weight22(reg_weight2_14_2), .reg_activation12(reg_activation2_14_1), .reg_activation22(reg_activation2_14_2), .weight_en(weight_en));
SA22 U2_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_15_1), .partial_sum_in12(reg_psum1_15_2), .weight_in11(reg_weight1_15_1), .weight_in12(reg_weight1_15_2), .activation_in11(reg_activation2_14_1), .activation_in21(reg_activation2_14_2), .reg_partial_sum21(reg_psum2_15_1), .reg_partial_sum22(reg_psum2_15_2), .reg_weight21(reg_weight2_15_1), .reg_weight22(reg_weight2_15_2), .reg_activation12(reg_activation2_15_1), .reg_activation22(reg_activation2_15_2), .weight_en(weight_en));
SA22 U2_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_16_1), .partial_sum_in12(reg_psum1_16_2), .weight_in11(reg_weight1_16_1), .weight_in12(reg_weight1_16_2), .activation_in11(reg_activation2_15_1), .activation_in21(reg_activation2_15_2), .reg_partial_sum21(reg_psum2_16_1), .reg_partial_sum22(reg_psum2_16_2), .reg_weight21(reg_weight2_16_1), .reg_weight22(reg_weight2_16_2), .reg_activation12(reg_activation2_16_1), .reg_activation22(reg_activation2_16_2), .weight_en(weight_en));
SA22 U2_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_17_1), .partial_sum_in12(reg_psum1_17_2), .weight_in11(reg_weight1_17_1), .weight_in12(reg_weight1_17_2), .activation_in11(reg_activation2_16_1), .activation_in21(reg_activation2_16_2), .reg_partial_sum21(reg_psum2_17_1), .reg_partial_sum22(reg_psum2_17_2), .reg_weight21(reg_weight2_17_1), .reg_weight22(reg_weight2_17_2), .reg_activation12(reg_activation2_17_1), .reg_activation22(reg_activation2_17_2), .weight_en(weight_en));
SA22 U2_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_18_1), .partial_sum_in12(reg_psum1_18_2), .weight_in11(reg_weight1_18_1), .weight_in12(reg_weight1_18_2), .activation_in11(reg_activation2_17_1), .activation_in21(reg_activation2_17_2), .reg_partial_sum21(reg_psum2_18_1), .reg_partial_sum22(reg_psum2_18_2), .reg_weight21(reg_weight2_18_1), .reg_weight22(reg_weight2_18_2), .reg_activation12(reg_activation2_18_1), .reg_activation22(reg_activation2_18_2), .weight_en(weight_en));
SA22 U2_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_19_1), .partial_sum_in12(reg_psum1_19_2), .weight_in11(reg_weight1_19_1), .weight_in12(reg_weight1_19_2), .activation_in11(reg_activation2_18_1), .activation_in21(reg_activation2_18_2), .reg_partial_sum21(reg_psum2_19_1), .reg_partial_sum22(reg_psum2_19_2), .reg_weight21(reg_weight2_19_1), .reg_weight22(reg_weight2_19_2), .reg_activation12(reg_activation2_19_1), .reg_activation22(reg_activation2_19_2), .weight_en(weight_en));
SA22 U2_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_20_1), .partial_sum_in12(reg_psum1_20_2), .weight_in11(reg_weight1_20_1), .weight_in12(reg_weight1_20_2), .activation_in11(reg_activation2_19_1), .activation_in21(reg_activation2_19_2), .reg_partial_sum21(reg_psum2_20_1), .reg_partial_sum22(reg_psum2_20_2), .reg_weight21(reg_weight2_20_1), .reg_weight22(reg_weight2_20_2), .reg_activation12(reg_activation2_20_1), .reg_activation22(reg_activation2_20_2), .weight_en(weight_en));
SA22 U2_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_21_1), .partial_sum_in12(reg_psum1_21_2), .weight_in11(reg_weight1_21_1), .weight_in12(reg_weight1_21_2), .activation_in11(reg_activation2_20_1), .activation_in21(reg_activation2_20_2), .reg_partial_sum21(reg_psum2_21_1), .reg_partial_sum22(reg_psum2_21_2), .reg_weight21(reg_weight2_21_1), .reg_weight22(reg_weight2_21_2), .reg_activation12(reg_activation2_21_1), .reg_activation22(reg_activation2_21_2), .weight_en(weight_en));
SA22 U2_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_22_1), .partial_sum_in12(reg_psum1_22_2), .weight_in11(reg_weight1_22_1), .weight_in12(reg_weight1_22_2), .activation_in11(reg_activation2_21_1), .activation_in21(reg_activation2_21_2), .reg_partial_sum21(reg_psum2_22_1), .reg_partial_sum22(reg_psum2_22_2), .reg_weight21(reg_weight2_22_1), .reg_weight22(reg_weight2_22_2), .reg_activation12(reg_activation2_22_1), .reg_activation22(reg_activation2_22_2), .weight_en(weight_en));
SA22 U2_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_23_1), .partial_sum_in12(reg_psum1_23_2), .weight_in11(reg_weight1_23_1), .weight_in12(reg_weight1_23_2), .activation_in11(reg_activation2_22_1), .activation_in21(reg_activation2_22_2), .reg_partial_sum21(reg_psum2_23_1), .reg_partial_sum22(reg_psum2_23_2), .reg_weight21(reg_weight2_23_1), .reg_weight22(reg_weight2_23_2), .reg_activation12(reg_activation2_23_1), .reg_activation22(reg_activation2_23_2), .weight_en(weight_en));
SA22 U2_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_24_1), .partial_sum_in12(reg_psum1_24_2), .weight_in11(reg_weight1_24_1), .weight_in12(reg_weight1_24_2), .activation_in11(reg_activation2_23_1), .activation_in21(reg_activation2_23_2), .reg_partial_sum21(reg_psum2_24_1), .reg_partial_sum22(reg_psum2_24_2), .reg_weight21(reg_weight2_24_1), .reg_weight22(reg_weight2_24_2), .reg_activation12(reg_activation2_24_1), .reg_activation22(reg_activation2_24_2), .weight_en(weight_en));
SA22 U2_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_25_1), .partial_sum_in12(reg_psum1_25_2), .weight_in11(reg_weight1_25_1), .weight_in12(reg_weight1_25_2), .activation_in11(reg_activation2_24_1), .activation_in21(reg_activation2_24_2), .reg_partial_sum21(reg_psum2_25_1), .reg_partial_sum22(reg_psum2_25_2), .reg_weight21(reg_weight2_25_1), .reg_weight22(reg_weight2_25_2), .reg_activation12(reg_activation2_25_1), .reg_activation22(reg_activation2_25_2), .weight_en(weight_en));
SA22 U2_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_26_1), .partial_sum_in12(reg_psum1_26_2), .weight_in11(reg_weight1_26_1), .weight_in12(reg_weight1_26_2), .activation_in11(reg_activation2_25_1), .activation_in21(reg_activation2_25_2), .reg_partial_sum21(reg_psum2_26_1), .reg_partial_sum22(reg_psum2_26_2), .reg_weight21(reg_weight2_26_1), .reg_weight22(reg_weight2_26_2), .reg_activation12(reg_activation2_26_1), .reg_activation22(reg_activation2_26_2), .weight_en(weight_en));
SA22 U2_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_27_1), .partial_sum_in12(reg_psum1_27_2), .weight_in11(reg_weight1_27_1), .weight_in12(reg_weight1_27_2), .activation_in11(reg_activation2_26_1), .activation_in21(reg_activation2_26_2), .reg_partial_sum21(reg_psum2_27_1), .reg_partial_sum22(reg_psum2_27_2), .reg_weight21(reg_weight2_27_1), .reg_weight22(reg_weight2_27_2), .reg_activation12(reg_activation2_27_1), .reg_activation22(reg_activation2_27_2), .weight_en(weight_en));
SA22 U2_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_28_1), .partial_sum_in12(reg_psum1_28_2), .weight_in11(reg_weight1_28_1), .weight_in12(reg_weight1_28_2), .activation_in11(reg_activation2_27_1), .activation_in21(reg_activation2_27_2), .reg_partial_sum21(reg_psum2_28_1), .reg_partial_sum22(reg_psum2_28_2), .reg_weight21(reg_weight2_28_1), .reg_weight22(reg_weight2_28_2), .reg_activation12(reg_activation2_28_1), .reg_activation22(reg_activation2_28_2), .weight_en(weight_en));
SA22 U2_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_29_1), .partial_sum_in12(reg_psum1_29_2), .weight_in11(reg_weight1_29_1), .weight_in12(reg_weight1_29_2), .activation_in11(reg_activation2_28_1), .activation_in21(reg_activation2_28_2), .reg_partial_sum21(reg_psum2_29_1), .reg_partial_sum22(reg_psum2_29_2), .reg_weight21(reg_weight2_29_1), .reg_weight22(reg_weight2_29_2), .reg_activation12(reg_activation2_29_1), .reg_activation22(reg_activation2_29_2), .weight_en(weight_en));
SA22 U2_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_30_1), .partial_sum_in12(reg_psum1_30_2), .weight_in11(reg_weight1_30_1), .weight_in12(reg_weight1_30_2), .activation_in11(reg_activation2_29_1), .activation_in21(reg_activation2_29_2), .reg_partial_sum21(reg_psum2_30_1), .reg_partial_sum22(reg_psum2_30_2), .reg_weight21(reg_weight2_30_1), .reg_weight22(reg_weight2_30_2), .reg_activation12(reg_activation2_30_1), .reg_activation22(reg_activation2_30_2), .weight_en(weight_en));
SA22 U2_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_31_1), .partial_sum_in12(reg_psum1_31_2), .weight_in11(reg_weight1_31_1), .weight_in12(reg_weight1_31_2), .activation_in11(reg_activation2_30_1), .activation_in21(reg_activation2_30_2), .reg_partial_sum21(reg_psum2_31_1), .reg_partial_sum22(reg_psum2_31_2), .reg_weight21(reg_weight2_31_1), .reg_weight22(reg_weight2_31_2), .reg_activation12(reg_activation2_31_1), .reg_activation22(reg_activation2_31_2), .weight_en(weight_en));
SA22 U2_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum1_32_1), .partial_sum_in12(reg_psum1_32_2), .weight_in11(reg_weight1_32_1), .weight_in12(reg_weight1_32_2), .activation_in11(reg_activation2_31_1), .activation_in21(reg_activation2_31_2), .reg_partial_sum21(reg_psum2_32_1), .reg_partial_sum22(reg_psum2_32_2), .reg_weight21(reg_weight2_32_1), .reg_weight22(reg_weight2_32_2), .weight_en(weight_en));
SA22 U3_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_1_1), .partial_sum_in12(reg_psum2_1_2), .weight_in11(reg_weight2_1_1), .weight_in12(reg_weight2_1_2), .activation_in11(in_activation3_1_1), .activation_in21(in_activation3_1_2), .reg_partial_sum21(reg_psum3_1_1), .reg_partial_sum22(reg_psum3_1_2), .reg_weight21(reg_weight3_1_1), .reg_weight22(reg_weight3_1_2), .reg_activation12(reg_activation3_1_1), .reg_activation22(reg_activation3_1_2), .weight_en(weight_en));
SA22 U3_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_2_1), .partial_sum_in12(reg_psum2_2_2), .weight_in11(reg_weight2_2_1), .weight_in12(reg_weight2_2_2), .activation_in11(reg_activation3_1_1), .activation_in21(reg_activation3_1_2), .reg_partial_sum21(reg_psum3_2_1), .reg_partial_sum22(reg_psum3_2_2), .reg_weight21(reg_weight3_2_1), .reg_weight22(reg_weight3_2_2), .reg_activation12(reg_activation3_2_1), .reg_activation22(reg_activation3_2_2), .weight_en(weight_en));
SA22 U3_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_3_1), .partial_sum_in12(reg_psum2_3_2), .weight_in11(reg_weight2_3_1), .weight_in12(reg_weight2_3_2), .activation_in11(reg_activation3_2_1), .activation_in21(reg_activation3_2_2), .reg_partial_sum21(reg_psum3_3_1), .reg_partial_sum22(reg_psum3_3_2), .reg_weight21(reg_weight3_3_1), .reg_weight22(reg_weight3_3_2), .reg_activation12(reg_activation3_3_1), .reg_activation22(reg_activation3_3_2), .weight_en(weight_en));
SA22 U3_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_4_1), .partial_sum_in12(reg_psum2_4_2), .weight_in11(reg_weight2_4_1), .weight_in12(reg_weight2_4_2), .activation_in11(reg_activation3_3_1), .activation_in21(reg_activation3_3_2), .reg_partial_sum21(reg_psum3_4_1), .reg_partial_sum22(reg_psum3_4_2), .reg_weight21(reg_weight3_4_1), .reg_weight22(reg_weight3_4_2), .reg_activation12(reg_activation3_4_1), .reg_activation22(reg_activation3_4_2), .weight_en(weight_en));
SA22 U3_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_5_1), .partial_sum_in12(reg_psum2_5_2), .weight_in11(reg_weight2_5_1), .weight_in12(reg_weight2_5_2), .activation_in11(reg_activation3_4_1), .activation_in21(reg_activation3_4_2), .reg_partial_sum21(reg_psum3_5_1), .reg_partial_sum22(reg_psum3_5_2), .reg_weight21(reg_weight3_5_1), .reg_weight22(reg_weight3_5_2), .reg_activation12(reg_activation3_5_1), .reg_activation22(reg_activation3_5_2), .weight_en(weight_en));
SA22 U3_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_6_1), .partial_sum_in12(reg_psum2_6_2), .weight_in11(reg_weight2_6_1), .weight_in12(reg_weight2_6_2), .activation_in11(reg_activation3_5_1), .activation_in21(reg_activation3_5_2), .reg_partial_sum21(reg_psum3_6_1), .reg_partial_sum22(reg_psum3_6_2), .reg_weight21(reg_weight3_6_1), .reg_weight22(reg_weight3_6_2), .reg_activation12(reg_activation3_6_1), .reg_activation22(reg_activation3_6_2), .weight_en(weight_en));
SA22 U3_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_7_1), .partial_sum_in12(reg_psum2_7_2), .weight_in11(reg_weight2_7_1), .weight_in12(reg_weight2_7_2), .activation_in11(reg_activation3_6_1), .activation_in21(reg_activation3_6_2), .reg_partial_sum21(reg_psum3_7_1), .reg_partial_sum22(reg_psum3_7_2), .reg_weight21(reg_weight3_7_1), .reg_weight22(reg_weight3_7_2), .reg_activation12(reg_activation3_7_1), .reg_activation22(reg_activation3_7_2), .weight_en(weight_en));
SA22 U3_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_8_1), .partial_sum_in12(reg_psum2_8_2), .weight_in11(reg_weight2_8_1), .weight_in12(reg_weight2_8_2), .activation_in11(reg_activation3_7_1), .activation_in21(reg_activation3_7_2), .reg_partial_sum21(reg_psum3_8_1), .reg_partial_sum22(reg_psum3_8_2), .reg_weight21(reg_weight3_8_1), .reg_weight22(reg_weight3_8_2), .reg_activation12(reg_activation3_8_1), .reg_activation22(reg_activation3_8_2), .weight_en(weight_en));
SA22 U3_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_9_1), .partial_sum_in12(reg_psum2_9_2), .weight_in11(reg_weight2_9_1), .weight_in12(reg_weight2_9_2), .activation_in11(reg_activation3_8_1), .activation_in21(reg_activation3_8_2), .reg_partial_sum21(reg_psum3_9_1), .reg_partial_sum22(reg_psum3_9_2), .reg_weight21(reg_weight3_9_1), .reg_weight22(reg_weight3_9_2), .reg_activation12(reg_activation3_9_1), .reg_activation22(reg_activation3_9_2), .weight_en(weight_en));
SA22 U3_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_10_1), .partial_sum_in12(reg_psum2_10_2), .weight_in11(reg_weight2_10_1), .weight_in12(reg_weight2_10_2), .activation_in11(reg_activation3_9_1), .activation_in21(reg_activation3_9_2), .reg_partial_sum21(reg_psum3_10_1), .reg_partial_sum22(reg_psum3_10_2), .reg_weight21(reg_weight3_10_1), .reg_weight22(reg_weight3_10_2), .reg_activation12(reg_activation3_10_1), .reg_activation22(reg_activation3_10_2), .weight_en(weight_en));
SA22 U3_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_11_1), .partial_sum_in12(reg_psum2_11_2), .weight_in11(reg_weight2_11_1), .weight_in12(reg_weight2_11_2), .activation_in11(reg_activation3_10_1), .activation_in21(reg_activation3_10_2), .reg_partial_sum21(reg_psum3_11_1), .reg_partial_sum22(reg_psum3_11_2), .reg_weight21(reg_weight3_11_1), .reg_weight22(reg_weight3_11_2), .reg_activation12(reg_activation3_11_1), .reg_activation22(reg_activation3_11_2), .weight_en(weight_en));
SA22 U3_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_12_1), .partial_sum_in12(reg_psum2_12_2), .weight_in11(reg_weight2_12_1), .weight_in12(reg_weight2_12_2), .activation_in11(reg_activation3_11_1), .activation_in21(reg_activation3_11_2), .reg_partial_sum21(reg_psum3_12_1), .reg_partial_sum22(reg_psum3_12_2), .reg_weight21(reg_weight3_12_1), .reg_weight22(reg_weight3_12_2), .reg_activation12(reg_activation3_12_1), .reg_activation22(reg_activation3_12_2), .weight_en(weight_en));
SA22 U3_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_13_1), .partial_sum_in12(reg_psum2_13_2), .weight_in11(reg_weight2_13_1), .weight_in12(reg_weight2_13_2), .activation_in11(reg_activation3_12_1), .activation_in21(reg_activation3_12_2), .reg_partial_sum21(reg_psum3_13_1), .reg_partial_sum22(reg_psum3_13_2), .reg_weight21(reg_weight3_13_1), .reg_weight22(reg_weight3_13_2), .reg_activation12(reg_activation3_13_1), .reg_activation22(reg_activation3_13_2), .weight_en(weight_en));
SA22 U3_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_14_1), .partial_sum_in12(reg_psum2_14_2), .weight_in11(reg_weight2_14_1), .weight_in12(reg_weight2_14_2), .activation_in11(reg_activation3_13_1), .activation_in21(reg_activation3_13_2), .reg_partial_sum21(reg_psum3_14_1), .reg_partial_sum22(reg_psum3_14_2), .reg_weight21(reg_weight3_14_1), .reg_weight22(reg_weight3_14_2), .reg_activation12(reg_activation3_14_1), .reg_activation22(reg_activation3_14_2), .weight_en(weight_en));
SA22 U3_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_15_1), .partial_sum_in12(reg_psum2_15_2), .weight_in11(reg_weight2_15_1), .weight_in12(reg_weight2_15_2), .activation_in11(reg_activation3_14_1), .activation_in21(reg_activation3_14_2), .reg_partial_sum21(reg_psum3_15_1), .reg_partial_sum22(reg_psum3_15_2), .reg_weight21(reg_weight3_15_1), .reg_weight22(reg_weight3_15_2), .reg_activation12(reg_activation3_15_1), .reg_activation22(reg_activation3_15_2), .weight_en(weight_en));
SA22 U3_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_16_1), .partial_sum_in12(reg_psum2_16_2), .weight_in11(reg_weight2_16_1), .weight_in12(reg_weight2_16_2), .activation_in11(reg_activation3_15_1), .activation_in21(reg_activation3_15_2), .reg_partial_sum21(reg_psum3_16_1), .reg_partial_sum22(reg_psum3_16_2), .reg_weight21(reg_weight3_16_1), .reg_weight22(reg_weight3_16_2), .reg_activation12(reg_activation3_16_1), .reg_activation22(reg_activation3_16_2), .weight_en(weight_en));
SA22 U3_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_17_1), .partial_sum_in12(reg_psum2_17_2), .weight_in11(reg_weight2_17_1), .weight_in12(reg_weight2_17_2), .activation_in11(reg_activation3_16_1), .activation_in21(reg_activation3_16_2), .reg_partial_sum21(reg_psum3_17_1), .reg_partial_sum22(reg_psum3_17_2), .reg_weight21(reg_weight3_17_1), .reg_weight22(reg_weight3_17_2), .reg_activation12(reg_activation3_17_1), .reg_activation22(reg_activation3_17_2), .weight_en(weight_en));
SA22 U3_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_18_1), .partial_sum_in12(reg_psum2_18_2), .weight_in11(reg_weight2_18_1), .weight_in12(reg_weight2_18_2), .activation_in11(reg_activation3_17_1), .activation_in21(reg_activation3_17_2), .reg_partial_sum21(reg_psum3_18_1), .reg_partial_sum22(reg_psum3_18_2), .reg_weight21(reg_weight3_18_1), .reg_weight22(reg_weight3_18_2), .reg_activation12(reg_activation3_18_1), .reg_activation22(reg_activation3_18_2), .weight_en(weight_en));
SA22 U3_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_19_1), .partial_sum_in12(reg_psum2_19_2), .weight_in11(reg_weight2_19_1), .weight_in12(reg_weight2_19_2), .activation_in11(reg_activation3_18_1), .activation_in21(reg_activation3_18_2), .reg_partial_sum21(reg_psum3_19_1), .reg_partial_sum22(reg_psum3_19_2), .reg_weight21(reg_weight3_19_1), .reg_weight22(reg_weight3_19_2), .reg_activation12(reg_activation3_19_1), .reg_activation22(reg_activation3_19_2), .weight_en(weight_en));
SA22 U3_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_20_1), .partial_sum_in12(reg_psum2_20_2), .weight_in11(reg_weight2_20_1), .weight_in12(reg_weight2_20_2), .activation_in11(reg_activation3_19_1), .activation_in21(reg_activation3_19_2), .reg_partial_sum21(reg_psum3_20_1), .reg_partial_sum22(reg_psum3_20_2), .reg_weight21(reg_weight3_20_1), .reg_weight22(reg_weight3_20_2), .reg_activation12(reg_activation3_20_1), .reg_activation22(reg_activation3_20_2), .weight_en(weight_en));
SA22 U3_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_21_1), .partial_sum_in12(reg_psum2_21_2), .weight_in11(reg_weight2_21_1), .weight_in12(reg_weight2_21_2), .activation_in11(reg_activation3_20_1), .activation_in21(reg_activation3_20_2), .reg_partial_sum21(reg_psum3_21_1), .reg_partial_sum22(reg_psum3_21_2), .reg_weight21(reg_weight3_21_1), .reg_weight22(reg_weight3_21_2), .reg_activation12(reg_activation3_21_1), .reg_activation22(reg_activation3_21_2), .weight_en(weight_en));
SA22 U3_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_22_1), .partial_sum_in12(reg_psum2_22_2), .weight_in11(reg_weight2_22_1), .weight_in12(reg_weight2_22_2), .activation_in11(reg_activation3_21_1), .activation_in21(reg_activation3_21_2), .reg_partial_sum21(reg_psum3_22_1), .reg_partial_sum22(reg_psum3_22_2), .reg_weight21(reg_weight3_22_1), .reg_weight22(reg_weight3_22_2), .reg_activation12(reg_activation3_22_1), .reg_activation22(reg_activation3_22_2), .weight_en(weight_en));
SA22 U3_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_23_1), .partial_sum_in12(reg_psum2_23_2), .weight_in11(reg_weight2_23_1), .weight_in12(reg_weight2_23_2), .activation_in11(reg_activation3_22_1), .activation_in21(reg_activation3_22_2), .reg_partial_sum21(reg_psum3_23_1), .reg_partial_sum22(reg_psum3_23_2), .reg_weight21(reg_weight3_23_1), .reg_weight22(reg_weight3_23_2), .reg_activation12(reg_activation3_23_1), .reg_activation22(reg_activation3_23_2), .weight_en(weight_en));
SA22 U3_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_24_1), .partial_sum_in12(reg_psum2_24_2), .weight_in11(reg_weight2_24_1), .weight_in12(reg_weight2_24_2), .activation_in11(reg_activation3_23_1), .activation_in21(reg_activation3_23_2), .reg_partial_sum21(reg_psum3_24_1), .reg_partial_sum22(reg_psum3_24_2), .reg_weight21(reg_weight3_24_1), .reg_weight22(reg_weight3_24_2), .reg_activation12(reg_activation3_24_1), .reg_activation22(reg_activation3_24_2), .weight_en(weight_en));
SA22 U3_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_25_1), .partial_sum_in12(reg_psum2_25_2), .weight_in11(reg_weight2_25_1), .weight_in12(reg_weight2_25_2), .activation_in11(reg_activation3_24_1), .activation_in21(reg_activation3_24_2), .reg_partial_sum21(reg_psum3_25_1), .reg_partial_sum22(reg_psum3_25_2), .reg_weight21(reg_weight3_25_1), .reg_weight22(reg_weight3_25_2), .reg_activation12(reg_activation3_25_1), .reg_activation22(reg_activation3_25_2), .weight_en(weight_en));
SA22 U3_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_26_1), .partial_sum_in12(reg_psum2_26_2), .weight_in11(reg_weight2_26_1), .weight_in12(reg_weight2_26_2), .activation_in11(reg_activation3_25_1), .activation_in21(reg_activation3_25_2), .reg_partial_sum21(reg_psum3_26_1), .reg_partial_sum22(reg_psum3_26_2), .reg_weight21(reg_weight3_26_1), .reg_weight22(reg_weight3_26_2), .reg_activation12(reg_activation3_26_1), .reg_activation22(reg_activation3_26_2), .weight_en(weight_en));
SA22 U3_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_27_1), .partial_sum_in12(reg_psum2_27_2), .weight_in11(reg_weight2_27_1), .weight_in12(reg_weight2_27_2), .activation_in11(reg_activation3_26_1), .activation_in21(reg_activation3_26_2), .reg_partial_sum21(reg_psum3_27_1), .reg_partial_sum22(reg_psum3_27_2), .reg_weight21(reg_weight3_27_1), .reg_weight22(reg_weight3_27_2), .reg_activation12(reg_activation3_27_1), .reg_activation22(reg_activation3_27_2), .weight_en(weight_en));
SA22 U3_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_28_1), .partial_sum_in12(reg_psum2_28_2), .weight_in11(reg_weight2_28_1), .weight_in12(reg_weight2_28_2), .activation_in11(reg_activation3_27_1), .activation_in21(reg_activation3_27_2), .reg_partial_sum21(reg_psum3_28_1), .reg_partial_sum22(reg_psum3_28_2), .reg_weight21(reg_weight3_28_1), .reg_weight22(reg_weight3_28_2), .reg_activation12(reg_activation3_28_1), .reg_activation22(reg_activation3_28_2), .weight_en(weight_en));
SA22 U3_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_29_1), .partial_sum_in12(reg_psum2_29_2), .weight_in11(reg_weight2_29_1), .weight_in12(reg_weight2_29_2), .activation_in11(reg_activation3_28_1), .activation_in21(reg_activation3_28_2), .reg_partial_sum21(reg_psum3_29_1), .reg_partial_sum22(reg_psum3_29_2), .reg_weight21(reg_weight3_29_1), .reg_weight22(reg_weight3_29_2), .reg_activation12(reg_activation3_29_1), .reg_activation22(reg_activation3_29_2), .weight_en(weight_en));
SA22 U3_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_30_1), .partial_sum_in12(reg_psum2_30_2), .weight_in11(reg_weight2_30_1), .weight_in12(reg_weight2_30_2), .activation_in11(reg_activation3_29_1), .activation_in21(reg_activation3_29_2), .reg_partial_sum21(reg_psum3_30_1), .reg_partial_sum22(reg_psum3_30_2), .reg_weight21(reg_weight3_30_1), .reg_weight22(reg_weight3_30_2), .reg_activation12(reg_activation3_30_1), .reg_activation22(reg_activation3_30_2), .weight_en(weight_en));
SA22 U3_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_31_1), .partial_sum_in12(reg_psum2_31_2), .weight_in11(reg_weight2_31_1), .weight_in12(reg_weight2_31_2), .activation_in11(reg_activation3_30_1), .activation_in21(reg_activation3_30_2), .reg_partial_sum21(reg_psum3_31_1), .reg_partial_sum22(reg_psum3_31_2), .reg_weight21(reg_weight3_31_1), .reg_weight22(reg_weight3_31_2), .reg_activation12(reg_activation3_31_1), .reg_activation22(reg_activation3_31_2), .weight_en(weight_en));
SA22 U3_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum2_32_1), .partial_sum_in12(reg_psum2_32_2), .weight_in11(reg_weight2_32_1), .weight_in12(reg_weight2_32_2), .activation_in11(reg_activation3_31_1), .activation_in21(reg_activation3_31_2), .reg_partial_sum21(reg_psum3_32_1), .reg_partial_sum22(reg_psum3_32_2), .reg_weight21(reg_weight3_32_1), .reg_weight22(reg_weight3_32_2), .weight_en(weight_en));
SA22 U4_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_1_1), .partial_sum_in12(reg_psum3_1_2), .weight_in11(reg_weight3_1_1), .weight_in12(reg_weight3_1_2), .activation_in11(in_activation4_1_1), .activation_in21(in_activation4_1_2), .reg_partial_sum21(reg_psum4_1_1), .reg_partial_sum22(reg_psum4_1_2), .reg_weight21(reg_weight4_1_1), .reg_weight22(reg_weight4_1_2), .reg_activation12(reg_activation4_1_1), .reg_activation22(reg_activation4_1_2), .weight_en(weight_en));
SA22 U4_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_2_1), .partial_sum_in12(reg_psum3_2_2), .weight_in11(reg_weight3_2_1), .weight_in12(reg_weight3_2_2), .activation_in11(reg_activation4_1_1), .activation_in21(reg_activation4_1_2), .reg_partial_sum21(reg_psum4_2_1), .reg_partial_sum22(reg_psum4_2_2), .reg_weight21(reg_weight4_2_1), .reg_weight22(reg_weight4_2_2), .reg_activation12(reg_activation4_2_1), .reg_activation22(reg_activation4_2_2), .weight_en(weight_en));
SA22 U4_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_3_1), .partial_sum_in12(reg_psum3_3_2), .weight_in11(reg_weight3_3_1), .weight_in12(reg_weight3_3_2), .activation_in11(reg_activation4_2_1), .activation_in21(reg_activation4_2_2), .reg_partial_sum21(reg_psum4_3_1), .reg_partial_sum22(reg_psum4_3_2), .reg_weight21(reg_weight4_3_1), .reg_weight22(reg_weight4_3_2), .reg_activation12(reg_activation4_3_1), .reg_activation22(reg_activation4_3_2), .weight_en(weight_en));
SA22 U4_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_4_1), .partial_sum_in12(reg_psum3_4_2), .weight_in11(reg_weight3_4_1), .weight_in12(reg_weight3_4_2), .activation_in11(reg_activation4_3_1), .activation_in21(reg_activation4_3_2), .reg_partial_sum21(reg_psum4_4_1), .reg_partial_sum22(reg_psum4_4_2), .reg_weight21(reg_weight4_4_1), .reg_weight22(reg_weight4_4_2), .reg_activation12(reg_activation4_4_1), .reg_activation22(reg_activation4_4_2), .weight_en(weight_en));
SA22 U4_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_5_1), .partial_sum_in12(reg_psum3_5_2), .weight_in11(reg_weight3_5_1), .weight_in12(reg_weight3_5_2), .activation_in11(reg_activation4_4_1), .activation_in21(reg_activation4_4_2), .reg_partial_sum21(reg_psum4_5_1), .reg_partial_sum22(reg_psum4_5_2), .reg_weight21(reg_weight4_5_1), .reg_weight22(reg_weight4_5_2), .reg_activation12(reg_activation4_5_1), .reg_activation22(reg_activation4_5_2), .weight_en(weight_en));
SA22 U4_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_6_1), .partial_sum_in12(reg_psum3_6_2), .weight_in11(reg_weight3_6_1), .weight_in12(reg_weight3_6_2), .activation_in11(reg_activation4_5_1), .activation_in21(reg_activation4_5_2), .reg_partial_sum21(reg_psum4_6_1), .reg_partial_sum22(reg_psum4_6_2), .reg_weight21(reg_weight4_6_1), .reg_weight22(reg_weight4_6_2), .reg_activation12(reg_activation4_6_1), .reg_activation22(reg_activation4_6_2), .weight_en(weight_en));
SA22 U4_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_7_1), .partial_sum_in12(reg_psum3_7_2), .weight_in11(reg_weight3_7_1), .weight_in12(reg_weight3_7_2), .activation_in11(reg_activation4_6_1), .activation_in21(reg_activation4_6_2), .reg_partial_sum21(reg_psum4_7_1), .reg_partial_sum22(reg_psum4_7_2), .reg_weight21(reg_weight4_7_1), .reg_weight22(reg_weight4_7_2), .reg_activation12(reg_activation4_7_1), .reg_activation22(reg_activation4_7_2), .weight_en(weight_en));
SA22 U4_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_8_1), .partial_sum_in12(reg_psum3_8_2), .weight_in11(reg_weight3_8_1), .weight_in12(reg_weight3_8_2), .activation_in11(reg_activation4_7_1), .activation_in21(reg_activation4_7_2), .reg_partial_sum21(reg_psum4_8_1), .reg_partial_sum22(reg_psum4_8_2), .reg_weight21(reg_weight4_8_1), .reg_weight22(reg_weight4_8_2), .reg_activation12(reg_activation4_8_1), .reg_activation22(reg_activation4_8_2), .weight_en(weight_en));
SA22 U4_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_9_1), .partial_sum_in12(reg_psum3_9_2), .weight_in11(reg_weight3_9_1), .weight_in12(reg_weight3_9_2), .activation_in11(reg_activation4_8_1), .activation_in21(reg_activation4_8_2), .reg_partial_sum21(reg_psum4_9_1), .reg_partial_sum22(reg_psum4_9_2), .reg_weight21(reg_weight4_9_1), .reg_weight22(reg_weight4_9_2), .reg_activation12(reg_activation4_9_1), .reg_activation22(reg_activation4_9_2), .weight_en(weight_en));
SA22 U4_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_10_1), .partial_sum_in12(reg_psum3_10_2), .weight_in11(reg_weight3_10_1), .weight_in12(reg_weight3_10_2), .activation_in11(reg_activation4_9_1), .activation_in21(reg_activation4_9_2), .reg_partial_sum21(reg_psum4_10_1), .reg_partial_sum22(reg_psum4_10_2), .reg_weight21(reg_weight4_10_1), .reg_weight22(reg_weight4_10_2), .reg_activation12(reg_activation4_10_1), .reg_activation22(reg_activation4_10_2), .weight_en(weight_en));
SA22 U4_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_11_1), .partial_sum_in12(reg_psum3_11_2), .weight_in11(reg_weight3_11_1), .weight_in12(reg_weight3_11_2), .activation_in11(reg_activation4_10_1), .activation_in21(reg_activation4_10_2), .reg_partial_sum21(reg_psum4_11_1), .reg_partial_sum22(reg_psum4_11_2), .reg_weight21(reg_weight4_11_1), .reg_weight22(reg_weight4_11_2), .reg_activation12(reg_activation4_11_1), .reg_activation22(reg_activation4_11_2), .weight_en(weight_en));
SA22 U4_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_12_1), .partial_sum_in12(reg_psum3_12_2), .weight_in11(reg_weight3_12_1), .weight_in12(reg_weight3_12_2), .activation_in11(reg_activation4_11_1), .activation_in21(reg_activation4_11_2), .reg_partial_sum21(reg_psum4_12_1), .reg_partial_sum22(reg_psum4_12_2), .reg_weight21(reg_weight4_12_1), .reg_weight22(reg_weight4_12_2), .reg_activation12(reg_activation4_12_1), .reg_activation22(reg_activation4_12_2), .weight_en(weight_en));
SA22 U4_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_13_1), .partial_sum_in12(reg_psum3_13_2), .weight_in11(reg_weight3_13_1), .weight_in12(reg_weight3_13_2), .activation_in11(reg_activation4_12_1), .activation_in21(reg_activation4_12_2), .reg_partial_sum21(reg_psum4_13_1), .reg_partial_sum22(reg_psum4_13_2), .reg_weight21(reg_weight4_13_1), .reg_weight22(reg_weight4_13_2), .reg_activation12(reg_activation4_13_1), .reg_activation22(reg_activation4_13_2), .weight_en(weight_en));
SA22 U4_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_14_1), .partial_sum_in12(reg_psum3_14_2), .weight_in11(reg_weight3_14_1), .weight_in12(reg_weight3_14_2), .activation_in11(reg_activation4_13_1), .activation_in21(reg_activation4_13_2), .reg_partial_sum21(reg_psum4_14_1), .reg_partial_sum22(reg_psum4_14_2), .reg_weight21(reg_weight4_14_1), .reg_weight22(reg_weight4_14_2), .reg_activation12(reg_activation4_14_1), .reg_activation22(reg_activation4_14_2), .weight_en(weight_en));
SA22 U4_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_15_1), .partial_sum_in12(reg_psum3_15_2), .weight_in11(reg_weight3_15_1), .weight_in12(reg_weight3_15_2), .activation_in11(reg_activation4_14_1), .activation_in21(reg_activation4_14_2), .reg_partial_sum21(reg_psum4_15_1), .reg_partial_sum22(reg_psum4_15_2), .reg_weight21(reg_weight4_15_1), .reg_weight22(reg_weight4_15_2), .reg_activation12(reg_activation4_15_1), .reg_activation22(reg_activation4_15_2), .weight_en(weight_en));
SA22 U4_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_16_1), .partial_sum_in12(reg_psum3_16_2), .weight_in11(reg_weight3_16_1), .weight_in12(reg_weight3_16_2), .activation_in11(reg_activation4_15_1), .activation_in21(reg_activation4_15_2), .reg_partial_sum21(reg_psum4_16_1), .reg_partial_sum22(reg_psum4_16_2), .reg_weight21(reg_weight4_16_1), .reg_weight22(reg_weight4_16_2), .reg_activation12(reg_activation4_16_1), .reg_activation22(reg_activation4_16_2), .weight_en(weight_en));
SA22 U4_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_17_1), .partial_sum_in12(reg_psum3_17_2), .weight_in11(reg_weight3_17_1), .weight_in12(reg_weight3_17_2), .activation_in11(reg_activation4_16_1), .activation_in21(reg_activation4_16_2), .reg_partial_sum21(reg_psum4_17_1), .reg_partial_sum22(reg_psum4_17_2), .reg_weight21(reg_weight4_17_1), .reg_weight22(reg_weight4_17_2), .reg_activation12(reg_activation4_17_1), .reg_activation22(reg_activation4_17_2), .weight_en(weight_en));
SA22 U4_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_18_1), .partial_sum_in12(reg_psum3_18_2), .weight_in11(reg_weight3_18_1), .weight_in12(reg_weight3_18_2), .activation_in11(reg_activation4_17_1), .activation_in21(reg_activation4_17_2), .reg_partial_sum21(reg_psum4_18_1), .reg_partial_sum22(reg_psum4_18_2), .reg_weight21(reg_weight4_18_1), .reg_weight22(reg_weight4_18_2), .reg_activation12(reg_activation4_18_1), .reg_activation22(reg_activation4_18_2), .weight_en(weight_en));
SA22 U4_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_19_1), .partial_sum_in12(reg_psum3_19_2), .weight_in11(reg_weight3_19_1), .weight_in12(reg_weight3_19_2), .activation_in11(reg_activation4_18_1), .activation_in21(reg_activation4_18_2), .reg_partial_sum21(reg_psum4_19_1), .reg_partial_sum22(reg_psum4_19_2), .reg_weight21(reg_weight4_19_1), .reg_weight22(reg_weight4_19_2), .reg_activation12(reg_activation4_19_1), .reg_activation22(reg_activation4_19_2), .weight_en(weight_en));
SA22 U4_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_20_1), .partial_sum_in12(reg_psum3_20_2), .weight_in11(reg_weight3_20_1), .weight_in12(reg_weight3_20_2), .activation_in11(reg_activation4_19_1), .activation_in21(reg_activation4_19_2), .reg_partial_sum21(reg_psum4_20_1), .reg_partial_sum22(reg_psum4_20_2), .reg_weight21(reg_weight4_20_1), .reg_weight22(reg_weight4_20_2), .reg_activation12(reg_activation4_20_1), .reg_activation22(reg_activation4_20_2), .weight_en(weight_en));
SA22 U4_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_21_1), .partial_sum_in12(reg_psum3_21_2), .weight_in11(reg_weight3_21_1), .weight_in12(reg_weight3_21_2), .activation_in11(reg_activation4_20_1), .activation_in21(reg_activation4_20_2), .reg_partial_sum21(reg_psum4_21_1), .reg_partial_sum22(reg_psum4_21_2), .reg_weight21(reg_weight4_21_1), .reg_weight22(reg_weight4_21_2), .reg_activation12(reg_activation4_21_1), .reg_activation22(reg_activation4_21_2), .weight_en(weight_en));
SA22 U4_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_22_1), .partial_sum_in12(reg_psum3_22_2), .weight_in11(reg_weight3_22_1), .weight_in12(reg_weight3_22_2), .activation_in11(reg_activation4_21_1), .activation_in21(reg_activation4_21_2), .reg_partial_sum21(reg_psum4_22_1), .reg_partial_sum22(reg_psum4_22_2), .reg_weight21(reg_weight4_22_1), .reg_weight22(reg_weight4_22_2), .reg_activation12(reg_activation4_22_1), .reg_activation22(reg_activation4_22_2), .weight_en(weight_en));
SA22 U4_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_23_1), .partial_sum_in12(reg_psum3_23_2), .weight_in11(reg_weight3_23_1), .weight_in12(reg_weight3_23_2), .activation_in11(reg_activation4_22_1), .activation_in21(reg_activation4_22_2), .reg_partial_sum21(reg_psum4_23_1), .reg_partial_sum22(reg_psum4_23_2), .reg_weight21(reg_weight4_23_1), .reg_weight22(reg_weight4_23_2), .reg_activation12(reg_activation4_23_1), .reg_activation22(reg_activation4_23_2), .weight_en(weight_en));
SA22 U4_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_24_1), .partial_sum_in12(reg_psum3_24_2), .weight_in11(reg_weight3_24_1), .weight_in12(reg_weight3_24_2), .activation_in11(reg_activation4_23_1), .activation_in21(reg_activation4_23_2), .reg_partial_sum21(reg_psum4_24_1), .reg_partial_sum22(reg_psum4_24_2), .reg_weight21(reg_weight4_24_1), .reg_weight22(reg_weight4_24_2), .reg_activation12(reg_activation4_24_1), .reg_activation22(reg_activation4_24_2), .weight_en(weight_en));
SA22 U4_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_25_1), .partial_sum_in12(reg_psum3_25_2), .weight_in11(reg_weight3_25_1), .weight_in12(reg_weight3_25_2), .activation_in11(reg_activation4_24_1), .activation_in21(reg_activation4_24_2), .reg_partial_sum21(reg_psum4_25_1), .reg_partial_sum22(reg_psum4_25_2), .reg_weight21(reg_weight4_25_1), .reg_weight22(reg_weight4_25_2), .reg_activation12(reg_activation4_25_1), .reg_activation22(reg_activation4_25_2), .weight_en(weight_en));
SA22 U4_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_26_1), .partial_sum_in12(reg_psum3_26_2), .weight_in11(reg_weight3_26_1), .weight_in12(reg_weight3_26_2), .activation_in11(reg_activation4_25_1), .activation_in21(reg_activation4_25_2), .reg_partial_sum21(reg_psum4_26_1), .reg_partial_sum22(reg_psum4_26_2), .reg_weight21(reg_weight4_26_1), .reg_weight22(reg_weight4_26_2), .reg_activation12(reg_activation4_26_1), .reg_activation22(reg_activation4_26_2), .weight_en(weight_en));
SA22 U4_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_27_1), .partial_sum_in12(reg_psum3_27_2), .weight_in11(reg_weight3_27_1), .weight_in12(reg_weight3_27_2), .activation_in11(reg_activation4_26_1), .activation_in21(reg_activation4_26_2), .reg_partial_sum21(reg_psum4_27_1), .reg_partial_sum22(reg_psum4_27_2), .reg_weight21(reg_weight4_27_1), .reg_weight22(reg_weight4_27_2), .reg_activation12(reg_activation4_27_1), .reg_activation22(reg_activation4_27_2), .weight_en(weight_en));
SA22 U4_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_28_1), .partial_sum_in12(reg_psum3_28_2), .weight_in11(reg_weight3_28_1), .weight_in12(reg_weight3_28_2), .activation_in11(reg_activation4_27_1), .activation_in21(reg_activation4_27_2), .reg_partial_sum21(reg_psum4_28_1), .reg_partial_sum22(reg_psum4_28_2), .reg_weight21(reg_weight4_28_1), .reg_weight22(reg_weight4_28_2), .reg_activation12(reg_activation4_28_1), .reg_activation22(reg_activation4_28_2), .weight_en(weight_en));
SA22 U4_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_29_1), .partial_sum_in12(reg_psum3_29_2), .weight_in11(reg_weight3_29_1), .weight_in12(reg_weight3_29_2), .activation_in11(reg_activation4_28_1), .activation_in21(reg_activation4_28_2), .reg_partial_sum21(reg_psum4_29_1), .reg_partial_sum22(reg_psum4_29_2), .reg_weight21(reg_weight4_29_1), .reg_weight22(reg_weight4_29_2), .reg_activation12(reg_activation4_29_1), .reg_activation22(reg_activation4_29_2), .weight_en(weight_en));
SA22 U4_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_30_1), .partial_sum_in12(reg_psum3_30_2), .weight_in11(reg_weight3_30_1), .weight_in12(reg_weight3_30_2), .activation_in11(reg_activation4_29_1), .activation_in21(reg_activation4_29_2), .reg_partial_sum21(reg_psum4_30_1), .reg_partial_sum22(reg_psum4_30_2), .reg_weight21(reg_weight4_30_1), .reg_weight22(reg_weight4_30_2), .reg_activation12(reg_activation4_30_1), .reg_activation22(reg_activation4_30_2), .weight_en(weight_en));
SA22 U4_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_31_1), .partial_sum_in12(reg_psum3_31_2), .weight_in11(reg_weight3_31_1), .weight_in12(reg_weight3_31_2), .activation_in11(reg_activation4_30_1), .activation_in21(reg_activation4_30_2), .reg_partial_sum21(reg_psum4_31_1), .reg_partial_sum22(reg_psum4_31_2), .reg_weight21(reg_weight4_31_1), .reg_weight22(reg_weight4_31_2), .reg_activation12(reg_activation4_31_1), .reg_activation22(reg_activation4_31_2), .weight_en(weight_en));
SA22 U4_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum3_32_1), .partial_sum_in12(reg_psum3_32_2), .weight_in11(reg_weight3_32_1), .weight_in12(reg_weight3_32_2), .activation_in11(reg_activation4_31_1), .activation_in21(reg_activation4_31_2), .reg_partial_sum21(reg_psum4_32_1), .reg_partial_sum22(reg_psum4_32_2), .reg_weight21(reg_weight4_32_1), .reg_weight22(reg_weight4_32_2), .weight_en(weight_en));
SA22 U5_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_1_1), .partial_sum_in12(reg_psum4_1_2), .weight_in11(reg_weight4_1_1), .weight_in12(reg_weight4_1_2), .activation_in11(in_activation5_1_1), .activation_in21(in_activation5_1_2), .reg_partial_sum21(reg_psum5_1_1), .reg_partial_sum22(reg_psum5_1_2), .reg_weight21(reg_weight5_1_1), .reg_weight22(reg_weight5_1_2), .reg_activation12(reg_activation5_1_1), .reg_activation22(reg_activation5_1_2), .weight_en(weight_en));
SA22 U5_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_2_1), .partial_sum_in12(reg_psum4_2_2), .weight_in11(reg_weight4_2_1), .weight_in12(reg_weight4_2_2), .activation_in11(reg_activation5_1_1), .activation_in21(reg_activation5_1_2), .reg_partial_sum21(reg_psum5_2_1), .reg_partial_sum22(reg_psum5_2_2), .reg_weight21(reg_weight5_2_1), .reg_weight22(reg_weight5_2_2), .reg_activation12(reg_activation5_2_1), .reg_activation22(reg_activation5_2_2), .weight_en(weight_en));
SA22 U5_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_3_1), .partial_sum_in12(reg_psum4_3_2), .weight_in11(reg_weight4_3_1), .weight_in12(reg_weight4_3_2), .activation_in11(reg_activation5_2_1), .activation_in21(reg_activation5_2_2), .reg_partial_sum21(reg_psum5_3_1), .reg_partial_sum22(reg_psum5_3_2), .reg_weight21(reg_weight5_3_1), .reg_weight22(reg_weight5_3_2), .reg_activation12(reg_activation5_3_1), .reg_activation22(reg_activation5_3_2), .weight_en(weight_en));
SA22 U5_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_4_1), .partial_sum_in12(reg_psum4_4_2), .weight_in11(reg_weight4_4_1), .weight_in12(reg_weight4_4_2), .activation_in11(reg_activation5_3_1), .activation_in21(reg_activation5_3_2), .reg_partial_sum21(reg_psum5_4_1), .reg_partial_sum22(reg_psum5_4_2), .reg_weight21(reg_weight5_4_1), .reg_weight22(reg_weight5_4_2), .reg_activation12(reg_activation5_4_1), .reg_activation22(reg_activation5_4_2), .weight_en(weight_en));
SA22 U5_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_5_1), .partial_sum_in12(reg_psum4_5_2), .weight_in11(reg_weight4_5_1), .weight_in12(reg_weight4_5_2), .activation_in11(reg_activation5_4_1), .activation_in21(reg_activation5_4_2), .reg_partial_sum21(reg_psum5_5_1), .reg_partial_sum22(reg_psum5_5_2), .reg_weight21(reg_weight5_5_1), .reg_weight22(reg_weight5_5_2), .reg_activation12(reg_activation5_5_1), .reg_activation22(reg_activation5_5_2), .weight_en(weight_en));
SA22 U5_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_6_1), .partial_sum_in12(reg_psum4_6_2), .weight_in11(reg_weight4_6_1), .weight_in12(reg_weight4_6_2), .activation_in11(reg_activation5_5_1), .activation_in21(reg_activation5_5_2), .reg_partial_sum21(reg_psum5_6_1), .reg_partial_sum22(reg_psum5_6_2), .reg_weight21(reg_weight5_6_1), .reg_weight22(reg_weight5_6_2), .reg_activation12(reg_activation5_6_1), .reg_activation22(reg_activation5_6_2), .weight_en(weight_en));
SA22 U5_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_7_1), .partial_sum_in12(reg_psum4_7_2), .weight_in11(reg_weight4_7_1), .weight_in12(reg_weight4_7_2), .activation_in11(reg_activation5_6_1), .activation_in21(reg_activation5_6_2), .reg_partial_sum21(reg_psum5_7_1), .reg_partial_sum22(reg_psum5_7_2), .reg_weight21(reg_weight5_7_1), .reg_weight22(reg_weight5_7_2), .reg_activation12(reg_activation5_7_1), .reg_activation22(reg_activation5_7_2), .weight_en(weight_en));
SA22 U5_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_8_1), .partial_sum_in12(reg_psum4_8_2), .weight_in11(reg_weight4_8_1), .weight_in12(reg_weight4_8_2), .activation_in11(reg_activation5_7_1), .activation_in21(reg_activation5_7_2), .reg_partial_sum21(reg_psum5_8_1), .reg_partial_sum22(reg_psum5_8_2), .reg_weight21(reg_weight5_8_1), .reg_weight22(reg_weight5_8_2), .reg_activation12(reg_activation5_8_1), .reg_activation22(reg_activation5_8_2), .weight_en(weight_en));
SA22 U5_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_9_1), .partial_sum_in12(reg_psum4_9_2), .weight_in11(reg_weight4_9_1), .weight_in12(reg_weight4_9_2), .activation_in11(reg_activation5_8_1), .activation_in21(reg_activation5_8_2), .reg_partial_sum21(reg_psum5_9_1), .reg_partial_sum22(reg_psum5_9_2), .reg_weight21(reg_weight5_9_1), .reg_weight22(reg_weight5_9_2), .reg_activation12(reg_activation5_9_1), .reg_activation22(reg_activation5_9_2), .weight_en(weight_en));
SA22 U5_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_10_1), .partial_sum_in12(reg_psum4_10_2), .weight_in11(reg_weight4_10_1), .weight_in12(reg_weight4_10_2), .activation_in11(reg_activation5_9_1), .activation_in21(reg_activation5_9_2), .reg_partial_sum21(reg_psum5_10_1), .reg_partial_sum22(reg_psum5_10_2), .reg_weight21(reg_weight5_10_1), .reg_weight22(reg_weight5_10_2), .reg_activation12(reg_activation5_10_1), .reg_activation22(reg_activation5_10_2), .weight_en(weight_en));
SA22 U5_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_11_1), .partial_sum_in12(reg_psum4_11_2), .weight_in11(reg_weight4_11_1), .weight_in12(reg_weight4_11_2), .activation_in11(reg_activation5_10_1), .activation_in21(reg_activation5_10_2), .reg_partial_sum21(reg_psum5_11_1), .reg_partial_sum22(reg_psum5_11_2), .reg_weight21(reg_weight5_11_1), .reg_weight22(reg_weight5_11_2), .reg_activation12(reg_activation5_11_1), .reg_activation22(reg_activation5_11_2), .weight_en(weight_en));
SA22 U5_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_12_1), .partial_sum_in12(reg_psum4_12_2), .weight_in11(reg_weight4_12_1), .weight_in12(reg_weight4_12_2), .activation_in11(reg_activation5_11_1), .activation_in21(reg_activation5_11_2), .reg_partial_sum21(reg_psum5_12_1), .reg_partial_sum22(reg_psum5_12_2), .reg_weight21(reg_weight5_12_1), .reg_weight22(reg_weight5_12_2), .reg_activation12(reg_activation5_12_1), .reg_activation22(reg_activation5_12_2), .weight_en(weight_en));
SA22 U5_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_13_1), .partial_sum_in12(reg_psum4_13_2), .weight_in11(reg_weight4_13_1), .weight_in12(reg_weight4_13_2), .activation_in11(reg_activation5_12_1), .activation_in21(reg_activation5_12_2), .reg_partial_sum21(reg_psum5_13_1), .reg_partial_sum22(reg_psum5_13_2), .reg_weight21(reg_weight5_13_1), .reg_weight22(reg_weight5_13_2), .reg_activation12(reg_activation5_13_1), .reg_activation22(reg_activation5_13_2), .weight_en(weight_en));
SA22 U5_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_14_1), .partial_sum_in12(reg_psum4_14_2), .weight_in11(reg_weight4_14_1), .weight_in12(reg_weight4_14_2), .activation_in11(reg_activation5_13_1), .activation_in21(reg_activation5_13_2), .reg_partial_sum21(reg_psum5_14_1), .reg_partial_sum22(reg_psum5_14_2), .reg_weight21(reg_weight5_14_1), .reg_weight22(reg_weight5_14_2), .reg_activation12(reg_activation5_14_1), .reg_activation22(reg_activation5_14_2), .weight_en(weight_en));
SA22 U5_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_15_1), .partial_sum_in12(reg_psum4_15_2), .weight_in11(reg_weight4_15_1), .weight_in12(reg_weight4_15_2), .activation_in11(reg_activation5_14_1), .activation_in21(reg_activation5_14_2), .reg_partial_sum21(reg_psum5_15_1), .reg_partial_sum22(reg_psum5_15_2), .reg_weight21(reg_weight5_15_1), .reg_weight22(reg_weight5_15_2), .reg_activation12(reg_activation5_15_1), .reg_activation22(reg_activation5_15_2), .weight_en(weight_en));
SA22 U5_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_16_1), .partial_sum_in12(reg_psum4_16_2), .weight_in11(reg_weight4_16_1), .weight_in12(reg_weight4_16_2), .activation_in11(reg_activation5_15_1), .activation_in21(reg_activation5_15_2), .reg_partial_sum21(reg_psum5_16_1), .reg_partial_sum22(reg_psum5_16_2), .reg_weight21(reg_weight5_16_1), .reg_weight22(reg_weight5_16_2), .reg_activation12(reg_activation5_16_1), .reg_activation22(reg_activation5_16_2), .weight_en(weight_en));
SA22 U5_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_17_1), .partial_sum_in12(reg_psum4_17_2), .weight_in11(reg_weight4_17_1), .weight_in12(reg_weight4_17_2), .activation_in11(reg_activation5_16_1), .activation_in21(reg_activation5_16_2), .reg_partial_sum21(reg_psum5_17_1), .reg_partial_sum22(reg_psum5_17_2), .reg_weight21(reg_weight5_17_1), .reg_weight22(reg_weight5_17_2), .reg_activation12(reg_activation5_17_1), .reg_activation22(reg_activation5_17_2), .weight_en(weight_en));
SA22 U5_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_18_1), .partial_sum_in12(reg_psum4_18_2), .weight_in11(reg_weight4_18_1), .weight_in12(reg_weight4_18_2), .activation_in11(reg_activation5_17_1), .activation_in21(reg_activation5_17_2), .reg_partial_sum21(reg_psum5_18_1), .reg_partial_sum22(reg_psum5_18_2), .reg_weight21(reg_weight5_18_1), .reg_weight22(reg_weight5_18_2), .reg_activation12(reg_activation5_18_1), .reg_activation22(reg_activation5_18_2), .weight_en(weight_en));
SA22 U5_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_19_1), .partial_sum_in12(reg_psum4_19_2), .weight_in11(reg_weight4_19_1), .weight_in12(reg_weight4_19_2), .activation_in11(reg_activation5_18_1), .activation_in21(reg_activation5_18_2), .reg_partial_sum21(reg_psum5_19_1), .reg_partial_sum22(reg_psum5_19_2), .reg_weight21(reg_weight5_19_1), .reg_weight22(reg_weight5_19_2), .reg_activation12(reg_activation5_19_1), .reg_activation22(reg_activation5_19_2), .weight_en(weight_en));
SA22 U5_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_20_1), .partial_sum_in12(reg_psum4_20_2), .weight_in11(reg_weight4_20_1), .weight_in12(reg_weight4_20_2), .activation_in11(reg_activation5_19_1), .activation_in21(reg_activation5_19_2), .reg_partial_sum21(reg_psum5_20_1), .reg_partial_sum22(reg_psum5_20_2), .reg_weight21(reg_weight5_20_1), .reg_weight22(reg_weight5_20_2), .reg_activation12(reg_activation5_20_1), .reg_activation22(reg_activation5_20_2), .weight_en(weight_en));
SA22 U5_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_21_1), .partial_sum_in12(reg_psum4_21_2), .weight_in11(reg_weight4_21_1), .weight_in12(reg_weight4_21_2), .activation_in11(reg_activation5_20_1), .activation_in21(reg_activation5_20_2), .reg_partial_sum21(reg_psum5_21_1), .reg_partial_sum22(reg_psum5_21_2), .reg_weight21(reg_weight5_21_1), .reg_weight22(reg_weight5_21_2), .reg_activation12(reg_activation5_21_1), .reg_activation22(reg_activation5_21_2), .weight_en(weight_en));
SA22 U5_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_22_1), .partial_sum_in12(reg_psum4_22_2), .weight_in11(reg_weight4_22_1), .weight_in12(reg_weight4_22_2), .activation_in11(reg_activation5_21_1), .activation_in21(reg_activation5_21_2), .reg_partial_sum21(reg_psum5_22_1), .reg_partial_sum22(reg_psum5_22_2), .reg_weight21(reg_weight5_22_1), .reg_weight22(reg_weight5_22_2), .reg_activation12(reg_activation5_22_1), .reg_activation22(reg_activation5_22_2), .weight_en(weight_en));
SA22 U5_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_23_1), .partial_sum_in12(reg_psum4_23_2), .weight_in11(reg_weight4_23_1), .weight_in12(reg_weight4_23_2), .activation_in11(reg_activation5_22_1), .activation_in21(reg_activation5_22_2), .reg_partial_sum21(reg_psum5_23_1), .reg_partial_sum22(reg_psum5_23_2), .reg_weight21(reg_weight5_23_1), .reg_weight22(reg_weight5_23_2), .reg_activation12(reg_activation5_23_1), .reg_activation22(reg_activation5_23_2), .weight_en(weight_en));
SA22 U5_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_24_1), .partial_sum_in12(reg_psum4_24_2), .weight_in11(reg_weight4_24_1), .weight_in12(reg_weight4_24_2), .activation_in11(reg_activation5_23_1), .activation_in21(reg_activation5_23_2), .reg_partial_sum21(reg_psum5_24_1), .reg_partial_sum22(reg_psum5_24_2), .reg_weight21(reg_weight5_24_1), .reg_weight22(reg_weight5_24_2), .reg_activation12(reg_activation5_24_1), .reg_activation22(reg_activation5_24_2), .weight_en(weight_en));
SA22 U5_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_25_1), .partial_sum_in12(reg_psum4_25_2), .weight_in11(reg_weight4_25_1), .weight_in12(reg_weight4_25_2), .activation_in11(reg_activation5_24_1), .activation_in21(reg_activation5_24_2), .reg_partial_sum21(reg_psum5_25_1), .reg_partial_sum22(reg_psum5_25_2), .reg_weight21(reg_weight5_25_1), .reg_weight22(reg_weight5_25_2), .reg_activation12(reg_activation5_25_1), .reg_activation22(reg_activation5_25_2), .weight_en(weight_en));
SA22 U5_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_26_1), .partial_sum_in12(reg_psum4_26_2), .weight_in11(reg_weight4_26_1), .weight_in12(reg_weight4_26_2), .activation_in11(reg_activation5_25_1), .activation_in21(reg_activation5_25_2), .reg_partial_sum21(reg_psum5_26_1), .reg_partial_sum22(reg_psum5_26_2), .reg_weight21(reg_weight5_26_1), .reg_weight22(reg_weight5_26_2), .reg_activation12(reg_activation5_26_1), .reg_activation22(reg_activation5_26_2), .weight_en(weight_en));
SA22 U5_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_27_1), .partial_sum_in12(reg_psum4_27_2), .weight_in11(reg_weight4_27_1), .weight_in12(reg_weight4_27_2), .activation_in11(reg_activation5_26_1), .activation_in21(reg_activation5_26_2), .reg_partial_sum21(reg_psum5_27_1), .reg_partial_sum22(reg_psum5_27_2), .reg_weight21(reg_weight5_27_1), .reg_weight22(reg_weight5_27_2), .reg_activation12(reg_activation5_27_1), .reg_activation22(reg_activation5_27_2), .weight_en(weight_en));
SA22 U5_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_28_1), .partial_sum_in12(reg_psum4_28_2), .weight_in11(reg_weight4_28_1), .weight_in12(reg_weight4_28_2), .activation_in11(reg_activation5_27_1), .activation_in21(reg_activation5_27_2), .reg_partial_sum21(reg_psum5_28_1), .reg_partial_sum22(reg_psum5_28_2), .reg_weight21(reg_weight5_28_1), .reg_weight22(reg_weight5_28_2), .reg_activation12(reg_activation5_28_1), .reg_activation22(reg_activation5_28_2), .weight_en(weight_en));
SA22 U5_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_29_1), .partial_sum_in12(reg_psum4_29_2), .weight_in11(reg_weight4_29_1), .weight_in12(reg_weight4_29_2), .activation_in11(reg_activation5_28_1), .activation_in21(reg_activation5_28_2), .reg_partial_sum21(reg_psum5_29_1), .reg_partial_sum22(reg_psum5_29_2), .reg_weight21(reg_weight5_29_1), .reg_weight22(reg_weight5_29_2), .reg_activation12(reg_activation5_29_1), .reg_activation22(reg_activation5_29_2), .weight_en(weight_en));
SA22 U5_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_30_1), .partial_sum_in12(reg_psum4_30_2), .weight_in11(reg_weight4_30_1), .weight_in12(reg_weight4_30_2), .activation_in11(reg_activation5_29_1), .activation_in21(reg_activation5_29_2), .reg_partial_sum21(reg_psum5_30_1), .reg_partial_sum22(reg_psum5_30_2), .reg_weight21(reg_weight5_30_1), .reg_weight22(reg_weight5_30_2), .reg_activation12(reg_activation5_30_1), .reg_activation22(reg_activation5_30_2), .weight_en(weight_en));
SA22 U5_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_31_1), .partial_sum_in12(reg_psum4_31_2), .weight_in11(reg_weight4_31_1), .weight_in12(reg_weight4_31_2), .activation_in11(reg_activation5_30_1), .activation_in21(reg_activation5_30_2), .reg_partial_sum21(reg_psum5_31_1), .reg_partial_sum22(reg_psum5_31_2), .reg_weight21(reg_weight5_31_1), .reg_weight22(reg_weight5_31_2), .reg_activation12(reg_activation5_31_1), .reg_activation22(reg_activation5_31_2), .weight_en(weight_en));
SA22 U5_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum4_32_1), .partial_sum_in12(reg_psum4_32_2), .weight_in11(reg_weight4_32_1), .weight_in12(reg_weight4_32_2), .activation_in11(reg_activation5_31_1), .activation_in21(reg_activation5_31_2), .reg_partial_sum21(reg_psum5_32_1), .reg_partial_sum22(reg_psum5_32_2), .reg_weight21(reg_weight5_32_1), .reg_weight22(reg_weight5_32_2), .weight_en(weight_en));
SA22 U6_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_1_1), .partial_sum_in12(reg_psum5_1_2), .weight_in11(reg_weight5_1_1), .weight_in12(reg_weight5_1_2), .activation_in11(in_activation6_1_1), .activation_in21(in_activation6_1_2), .reg_partial_sum21(reg_psum6_1_1), .reg_partial_sum22(reg_psum6_1_2), .reg_weight21(reg_weight6_1_1), .reg_weight22(reg_weight6_1_2), .reg_activation12(reg_activation6_1_1), .reg_activation22(reg_activation6_1_2), .weight_en(weight_en));
SA22 U6_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_2_1), .partial_sum_in12(reg_psum5_2_2), .weight_in11(reg_weight5_2_1), .weight_in12(reg_weight5_2_2), .activation_in11(reg_activation6_1_1), .activation_in21(reg_activation6_1_2), .reg_partial_sum21(reg_psum6_2_1), .reg_partial_sum22(reg_psum6_2_2), .reg_weight21(reg_weight6_2_1), .reg_weight22(reg_weight6_2_2), .reg_activation12(reg_activation6_2_1), .reg_activation22(reg_activation6_2_2), .weight_en(weight_en));
SA22 U6_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_3_1), .partial_sum_in12(reg_psum5_3_2), .weight_in11(reg_weight5_3_1), .weight_in12(reg_weight5_3_2), .activation_in11(reg_activation6_2_1), .activation_in21(reg_activation6_2_2), .reg_partial_sum21(reg_psum6_3_1), .reg_partial_sum22(reg_psum6_3_2), .reg_weight21(reg_weight6_3_1), .reg_weight22(reg_weight6_3_2), .reg_activation12(reg_activation6_3_1), .reg_activation22(reg_activation6_3_2), .weight_en(weight_en));
SA22 U6_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_4_1), .partial_sum_in12(reg_psum5_4_2), .weight_in11(reg_weight5_4_1), .weight_in12(reg_weight5_4_2), .activation_in11(reg_activation6_3_1), .activation_in21(reg_activation6_3_2), .reg_partial_sum21(reg_psum6_4_1), .reg_partial_sum22(reg_psum6_4_2), .reg_weight21(reg_weight6_4_1), .reg_weight22(reg_weight6_4_2), .reg_activation12(reg_activation6_4_1), .reg_activation22(reg_activation6_4_2), .weight_en(weight_en));
SA22 U6_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_5_1), .partial_sum_in12(reg_psum5_5_2), .weight_in11(reg_weight5_5_1), .weight_in12(reg_weight5_5_2), .activation_in11(reg_activation6_4_1), .activation_in21(reg_activation6_4_2), .reg_partial_sum21(reg_psum6_5_1), .reg_partial_sum22(reg_psum6_5_2), .reg_weight21(reg_weight6_5_1), .reg_weight22(reg_weight6_5_2), .reg_activation12(reg_activation6_5_1), .reg_activation22(reg_activation6_5_2), .weight_en(weight_en));
SA22 U6_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_6_1), .partial_sum_in12(reg_psum5_6_2), .weight_in11(reg_weight5_6_1), .weight_in12(reg_weight5_6_2), .activation_in11(reg_activation6_5_1), .activation_in21(reg_activation6_5_2), .reg_partial_sum21(reg_psum6_6_1), .reg_partial_sum22(reg_psum6_6_2), .reg_weight21(reg_weight6_6_1), .reg_weight22(reg_weight6_6_2), .reg_activation12(reg_activation6_6_1), .reg_activation22(reg_activation6_6_2), .weight_en(weight_en));
SA22 U6_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_7_1), .partial_sum_in12(reg_psum5_7_2), .weight_in11(reg_weight5_7_1), .weight_in12(reg_weight5_7_2), .activation_in11(reg_activation6_6_1), .activation_in21(reg_activation6_6_2), .reg_partial_sum21(reg_psum6_7_1), .reg_partial_sum22(reg_psum6_7_2), .reg_weight21(reg_weight6_7_1), .reg_weight22(reg_weight6_7_2), .reg_activation12(reg_activation6_7_1), .reg_activation22(reg_activation6_7_2), .weight_en(weight_en));
SA22 U6_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_8_1), .partial_sum_in12(reg_psum5_8_2), .weight_in11(reg_weight5_8_1), .weight_in12(reg_weight5_8_2), .activation_in11(reg_activation6_7_1), .activation_in21(reg_activation6_7_2), .reg_partial_sum21(reg_psum6_8_1), .reg_partial_sum22(reg_psum6_8_2), .reg_weight21(reg_weight6_8_1), .reg_weight22(reg_weight6_8_2), .reg_activation12(reg_activation6_8_1), .reg_activation22(reg_activation6_8_2), .weight_en(weight_en));
SA22 U6_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_9_1), .partial_sum_in12(reg_psum5_9_2), .weight_in11(reg_weight5_9_1), .weight_in12(reg_weight5_9_2), .activation_in11(reg_activation6_8_1), .activation_in21(reg_activation6_8_2), .reg_partial_sum21(reg_psum6_9_1), .reg_partial_sum22(reg_psum6_9_2), .reg_weight21(reg_weight6_9_1), .reg_weight22(reg_weight6_9_2), .reg_activation12(reg_activation6_9_1), .reg_activation22(reg_activation6_9_2), .weight_en(weight_en));
SA22 U6_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_10_1), .partial_sum_in12(reg_psum5_10_2), .weight_in11(reg_weight5_10_1), .weight_in12(reg_weight5_10_2), .activation_in11(reg_activation6_9_1), .activation_in21(reg_activation6_9_2), .reg_partial_sum21(reg_psum6_10_1), .reg_partial_sum22(reg_psum6_10_2), .reg_weight21(reg_weight6_10_1), .reg_weight22(reg_weight6_10_2), .reg_activation12(reg_activation6_10_1), .reg_activation22(reg_activation6_10_2), .weight_en(weight_en));
SA22 U6_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_11_1), .partial_sum_in12(reg_psum5_11_2), .weight_in11(reg_weight5_11_1), .weight_in12(reg_weight5_11_2), .activation_in11(reg_activation6_10_1), .activation_in21(reg_activation6_10_2), .reg_partial_sum21(reg_psum6_11_1), .reg_partial_sum22(reg_psum6_11_2), .reg_weight21(reg_weight6_11_1), .reg_weight22(reg_weight6_11_2), .reg_activation12(reg_activation6_11_1), .reg_activation22(reg_activation6_11_2), .weight_en(weight_en));
SA22 U6_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_12_1), .partial_sum_in12(reg_psum5_12_2), .weight_in11(reg_weight5_12_1), .weight_in12(reg_weight5_12_2), .activation_in11(reg_activation6_11_1), .activation_in21(reg_activation6_11_2), .reg_partial_sum21(reg_psum6_12_1), .reg_partial_sum22(reg_psum6_12_2), .reg_weight21(reg_weight6_12_1), .reg_weight22(reg_weight6_12_2), .reg_activation12(reg_activation6_12_1), .reg_activation22(reg_activation6_12_2), .weight_en(weight_en));
SA22 U6_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_13_1), .partial_sum_in12(reg_psum5_13_2), .weight_in11(reg_weight5_13_1), .weight_in12(reg_weight5_13_2), .activation_in11(reg_activation6_12_1), .activation_in21(reg_activation6_12_2), .reg_partial_sum21(reg_psum6_13_1), .reg_partial_sum22(reg_psum6_13_2), .reg_weight21(reg_weight6_13_1), .reg_weight22(reg_weight6_13_2), .reg_activation12(reg_activation6_13_1), .reg_activation22(reg_activation6_13_2), .weight_en(weight_en));
SA22 U6_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_14_1), .partial_sum_in12(reg_psum5_14_2), .weight_in11(reg_weight5_14_1), .weight_in12(reg_weight5_14_2), .activation_in11(reg_activation6_13_1), .activation_in21(reg_activation6_13_2), .reg_partial_sum21(reg_psum6_14_1), .reg_partial_sum22(reg_psum6_14_2), .reg_weight21(reg_weight6_14_1), .reg_weight22(reg_weight6_14_2), .reg_activation12(reg_activation6_14_1), .reg_activation22(reg_activation6_14_2), .weight_en(weight_en));
SA22 U6_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_15_1), .partial_sum_in12(reg_psum5_15_2), .weight_in11(reg_weight5_15_1), .weight_in12(reg_weight5_15_2), .activation_in11(reg_activation6_14_1), .activation_in21(reg_activation6_14_2), .reg_partial_sum21(reg_psum6_15_1), .reg_partial_sum22(reg_psum6_15_2), .reg_weight21(reg_weight6_15_1), .reg_weight22(reg_weight6_15_2), .reg_activation12(reg_activation6_15_1), .reg_activation22(reg_activation6_15_2), .weight_en(weight_en));
SA22 U6_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_16_1), .partial_sum_in12(reg_psum5_16_2), .weight_in11(reg_weight5_16_1), .weight_in12(reg_weight5_16_2), .activation_in11(reg_activation6_15_1), .activation_in21(reg_activation6_15_2), .reg_partial_sum21(reg_psum6_16_1), .reg_partial_sum22(reg_psum6_16_2), .reg_weight21(reg_weight6_16_1), .reg_weight22(reg_weight6_16_2), .reg_activation12(reg_activation6_16_1), .reg_activation22(reg_activation6_16_2), .weight_en(weight_en));
SA22 U6_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_17_1), .partial_sum_in12(reg_psum5_17_2), .weight_in11(reg_weight5_17_1), .weight_in12(reg_weight5_17_2), .activation_in11(reg_activation6_16_1), .activation_in21(reg_activation6_16_2), .reg_partial_sum21(reg_psum6_17_1), .reg_partial_sum22(reg_psum6_17_2), .reg_weight21(reg_weight6_17_1), .reg_weight22(reg_weight6_17_2), .reg_activation12(reg_activation6_17_1), .reg_activation22(reg_activation6_17_2), .weight_en(weight_en));
SA22 U6_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_18_1), .partial_sum_in12(reg_psum5_18_2), .weight_in11(reg_weight5_18_1), .weight_in12(reg_weight5_18_2), .activation_in11(reg_activation6_17_1), .activation_in21(reg_activation6_17_2), .reg_partial_sum21(reg_psum6_18_1), .reg_partial_sum22(reg_psum6_18_2), .reg_weight21(reg_weight6_18_1), .reg_weight22(reg_weight6_18_2), .reg_activation12(reg_activation6_18_1), .reg_activation22(reg_activation6_18_2), .weight_en(weight_en));
SA22 U6_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_19_1), .partial_sum_in12(reg_psum5_19_2), .weight_in11(reg_weight5_19_1), .weight_in12(reg_weight5_19_2), .activation_in11(reg_activation6_18_1), .activation_in21(reg_activation6_18_2), .reg_partial_sum21(reg_psum6_19_1), .reg_partial_sum22(reg_psum6_19_2), .reg_weight21(reg_weight6_19_1), .reg_weight22(reg_weight6_19_2), .reg_activation12(reg_activation6_19_1), .reg_activation22(reg_activation6_19_2), .weight_en(weight_en));
SA22 U6_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_20_1), .partial_sum_in12(reg_psum5_20_2), .weight_in11(reg_weight5_20_1), .weight_in12(reg_weight5_20_2), .activation_in11(reg_activation6_19_1), .activation_in21(reg_activation6_19_2), .reg_partial_sum21(reg_psum6_20_1), .reg_partial_sum22(reg_psum6_20_2), .reg_weight21(reg_weight6_20_1), .reg_weight22(reg_weight6_20_2), .reg_activation12(reg_activation6_20_1), .reg_activation22(reg_activation6_20_2), .weight_en(weight_en));
SA22 U6_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_21_1), .partial_sum_in12(reg_psum5_21_2), .weight_in11(reg_weight5_21_1), .weight_in12(reg_weight5_21_2), .activation_in11(reg_activation6_20_1), .activation_in21(reg_activation6_20_2), .reg_partial_sum21(reg_psum6_21_1), .reg_partial_sum22(reg_psum6_21_2), .reg_weight21(reg_weight6_21_1), .reg_weight22(reg_weight6_21_2), .reg_activation12(reg_activation6_21_1), .reg_activation22(reg_activation6_21_2), .weight_en(weight_en));
SA22 U6_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_22_1), .partial_sum_in12(reg_psum5_22_2), .weight_in11(reg_weight5_22_1), .weight_in12(reg_weight5_22_2), .activation_in11(reg_activation6_21_1), .activation_in21(reg_activation6_21_2), .reg_partial_sum21(reg_psum6_22_1), .reg_partial_sum22(reg_psum6_22_2), .reg_weight21(reg_weight6_22_1), .reg_weight22(reg_weight6_22_2), .reg_activation12(reg_activation6_22_1), .reg_activation22(reg_activation6_22_2), .weight_en(weight_en));
SA22 U6_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_23_1), .partial_sum_in12(reg_psum5_23_2), .weight_in11(reg_weight5_23_1), .weight_in12(reg_weight5_23_2), .activation_in11(reg_activation6_22_1), .activation_in21(reg_activation6_22_2), .reg_partial_sum21(reg_psum6_23_1), .reg_partial_sum22(reg_psum6_23_2), .reg_weight21(reg_weight6_23_1), .reg_weight22(reg_weight6_23_2), .reg_activation12(reg_activation6_23_1), .reg_activation22(reg_activation6_23_2), .weight_en(weight_en));
SA22 U6_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_24_1), .partial_sum_in12(reg_psum5_24_2), .weight_in11(reg_weight5_24_1), .weight_in12(reg_weight5_24_2), .activation_in11(reg_activation6_23_1), .activation_in21(reg_activation6_23_2), .reg_partial_sum21(reg_psum6_24_1), .reg_partial_sum22(reg_psum6_24_2), .reg_weight21(reg_weight6_24_1), .reg_weight22(reg_weight6_24_2), .reg_activation12(reg_activation6_24_1), .reg_activation22(reg_activation6_24_2), .weight_en(weight_en));
SA22 U6_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_25_1), .partial_sum_in12(reg_psum5_25_2), .weight_in11(reg_weight5_25_1), .weight_in12(reg_weight5_25_2), .activation_in11(reg_activation6_24_1), .activation_in21(reg_activation6_24_2), .reg_partial_sum21(reg_psum6_25_1), .reg_partial_sum22(reg_psum6_25_2), .reg_weight21(reg_weight6_25_1), .reg_weight22(reg_weight6_25_2), .reg_activation12(reg_activation6_25_1), .reg_activation22(reg_activation6_25_2), .weight_en(weight_en));
SA22 U6_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_26_1), .partial_sum_in12(reg_psum5_26_2), .weight_in11(reg_weight5_26_1), .weight_in12(reg_weight5_26_2), .activation_in11(reg_activation6_25_1), .activation_in21(reg_activation6_25_2), .reg_partial_sum21(reg_psum6_26_1), .reg_partial_sum22(reg_psum6_26_2), .reg_weight21(reg_weight6_26_1), .reg_weight22(reg_weight6_26_2), .reg_activation12(reg_activation6_26_1), .reg_activation22(reg_activation6_26_2), .weight_en(weight_en));
SA22 U6_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_27_1), .partial_sum_in12(reg_psum5_27_2), .weight_in11(reg_weight5_27_1), .weight_in12(reg_weight5_27_2), .activation_in11(reg_activation6_26_1), .activation_in21(reg_activation6_26_2), .reg_partial_sum21(reg_psum6_27_1), .reg_partial_sum22(reg_psum6_27_2), .reg_weight21(reg_weight6_27_1), .reg_weight22(reg_weight6_27_2), .reg_activation12(reg_activation6_27_1), .reg_activation22(reg_activation6_27_2), .weight_en(weight_en));
SA22 U6_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_28_1), .partial_sum_in12(reg_psum5_28_2), .weight_in11(reg_weight5_28_1), .weight_in12(reg_weight5_28_2), .activation_in11(reg_activation6_27_1), .activation_in21(reg_activation6_27_2), .reg_partial_sum21(reg_psum6_28_1), .reg_partial_sum22(reg_psum6_28_2), .reg_weight21(reg_weight6_28_1), .reg_weight22(reg_weight6_28_2), .reg_activation12(reg_activation6_28_1), .reg_activation22(reg_activation6_28_2), .weight_en(weight_en));
SA22 U6_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_29_1), .partial_sum_in12(reg_psum5_29_2), .weight_in11(reg_weight5_29_1), .weight_in12(reg_weight5_29_2), .activation_in11(reg_activation6_28_1), .activation_in21(reg_activation6_28_2), .reg_partial_sum21(reg_psum6_29_1), .reg_partial_sum22(reg_psum6_29_2), .reg_weight21(reg_weight6_29_1), .reg_weight22(reg_weight6_29_2), .reg_activation12(reg_activation6_29_1), .reg_activation22(reg_activation6_29_2), .weight_en(weight_en));
SA22 U6_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_30_1), .partial_sum_in12(reg_psum5_30_2), .weight_in11(reg_weight5_30_1), .weight_in12(reg_weight5_30_2), .activation_in11(reg_activation6_29_1), .activation_in21(reg_activation6_29_2), .reg_partial_sum21(reg_psum6_30_1), .reg_partial_sum22(reg_psum6_30_2), .reg_weight21(reg_weight6_30_1), .reg_weight22(reg_weight6_30_2), .reg_activation12(reg_activation6_30_1), .reg_activation22(reg_activation6_30_2), .weight_en(weight_en));
SA22 U6_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_31_1), .partial_sum_in12(reg_psum5_31_2), .weight_in11(reg_weight5_31_1), .weight_in12(reg_weight5_31_2), .activation_in11(reg_activation6_30_1), .activation_in21(reg_activation6_30_2), .reg_partial_sum21(reg_psum6_31_1), .reg_partial_sum22(reg_psum6_31_2), .reg_weight21(reg_weight6_31_1), .reg_weight22(reg_weight6_31_2), .reg_activation12(reg_activation6_31_1), .reg_activation22(reg_activation6_31_2), .weight_en(weight_en));
SA22 U6_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum5_32_1), .partial_sum_in12(reg_psum5_32_2), .weight_in11(reg_weight5_32_1), .weight_in12(reg_weight5_32_2), .activation_in11(reg_activation6_31_1), .activation_in21(reg_activation6_31_2), .reg_partial_sum21(reg_psum6_32_1), .reg_partial_sum22(reg_psum6_32_2), .reg_weight21(reg_weight6_32_1), .reg_weight22(reg_weight6_32_2), .weight_en(weight_en));
SA22 U7_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_1_1), .partial_sum_in12(reg_psum6_1_2), .weight_in11(reg_weight6_1_1), .weight_in12(reg_weight6_1_2), .activation_in11(in_activation7_1_1), .activation_in21(in_activation7_1_2), .reg_partial_sum21(reg_psum7_1_1), .reg_partial_sum22(reg_psum7_1_2), .reg_weight21(reg_weight7_1_1), .reg_weight22(reg_weight7_1_2), .reg_activation12(reg_activation7_1_1), .reg_activation22(reg_activation7_1_2), .weight_en(weight_en));
SA22 U7_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_2_1), .partial_sum_in12(reg_psum6_2_2), .weight_in11(reg_weight6_2_1), .weight_in12(reg_weight6_2_2), .activation_in11(reg_activation7_1_1), .activation_in21(reg_activation7_1_2), .reg_partial_sum21(reg_psum7_2_1), .reg_partial_sum22(reg_psum7_2_2), .reg_weight21(reg_weight7_2_1), .reg_weight22(reg_weight7_2_2), .reg_activation12(reg_activation7_2_1), .reg_activation22(reg_activation7_2_2), .weight_en(weight_en));
SA22 U7_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_3_1), .partial_sum_in12(reg_psum6_3_2), .weight_in11(reg_weight6_3_1), .weight_in12(reg_weight6_3_2), .activation_in11(reg_activation7_2_1), .activation_in21(reg_activation7_2_2), .reg_partial_sum21(reg_psum7_3_1), .reg_partial_sum22(reg_psum7_3_2), .reg_weight21(reg_weight7_3_1), .reg_weight22(reg_weight7_3_2), .reg_activation12(reg_activation7_3_1), .reg_activation22(reg_activation7_3_2), .weight_en(weight_en));
SA22 U7_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_4_1), .partial_sum_in12(reg_psum6_4_2), .weight_in11(reg_weight6_4_1), .weight_in12(reg_weight6_4_2), .activation_in11(reg_activation7_3_1), .activation_in21(reg_activation7_3_2), .reg_partial_sum21(reg_psum7_4_1), .reg_partial_sum22(reg_psum7_4_2), .reg_weight21(reg_weight7_4_1), .reg_weight22(reg_weight7_4_2), .reg_activation12(reg_activation7_4_1), .reg_activation22(reg_activation7_4_2), .weight_en(weight_en));
SA22 U7_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_5_1), .partial_sum_in12(reg_psum6_5_2), .weight_in11(reg_weight6_5_1), .weight_in12(reg_weight6_5_2), .activation_in11(reg_activation7_4_1), .activation_in21(reg_activation7_4_2), .reg_partial_sum21(reg_psum7_5_1), .reg_partial_sum22(reg_psum7_5_2), .reg_weight21(reg_weight7_5_1), .reg_weight22(reg_weight7_5_2), .reg_activation12(reg_activation7_5_1), .reg_activation22(reg_activation7_5_2), .weight_en(weight_en));
SA22 U7_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_6_1), .partial_sum_in12(reg_psum6_6_2), .weight_in11(reg_weight6_6_1), .weight_in12(reg_weight6_6_2), .activation_in11(reg_activation7_5_1), .activation_in21(reg_activation7_5_2), .reg_partial_sum21(reg_psum7_6_1), .reg_partial_sum22(reg_psum7_6_2), .reg_weight21(reg_weight7_6_1), .reg_weight22(reg_weight7_6_2), .reg_activation12(reg_activation7_6_1), .reg_activation22(reg_activation7_6_2), .weight_en(weight_en));
SA22 U7_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_7_1), .partial_sum_in12(reg_psum6_7_2), .weight_in11(reg_weight6_7_1), .weight_in12(reg_weight6_7_2), .activation_in11(reg_activation7_6_1), .activation_in21(reg_activation7_6_2), .reg_partial_sum21(reg_psum7_7_1), .reg_partial_sum22(reg_psum7_7_2), .reg_weight21(reg_weight7_7_1), .reg_weight22(reg_weight7_7_2), .reg_activation12(reg_activation7_7_1), .reg_activation22(reg_activation7_7_2), .weight_en(weight_en));
SA22 U7_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_8_1), .partial_sum_in12(reg_psum6_8_2), .weight_in11(reg_weight6_8_1), .weight_in12(reg_weight6_8_2), .activation_in11(reg_activation7_7_1), .activation_in21(reg_activation7_7_2), .reg_partial_sum21(reg_psum7_8_1), .reg_partial_sum22(reg_psum7_8_2), .reg_weight21(reg_weight7_8_1), .reg_weight22(reg_weight7_8_2), .reg_activation12(reg_activation7_8_1), .reg_activation22(reg_activation7_8_2), .weight_en(weight_en));
SA22 U7_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_9_1), .partial_sum_in12(reg_psum6_9_2), .weight_in11(reg_weight6_9_1), .weight_in12(reg_weight6_9_2), .activation_in11(reg_activation7_8_1), .activation_in21(reg_activation7_8_2), .reg_partial_sum21(reg_psum7_9_1), .reg_partial_sum22(reg_psum7_9_2), .reg_weight21(reg_weight7_9_1), .reg_weight22(reg_weight7_9_2), .reg_activation12(reg_activation7_9_1), .reg_activation22(reg_activation7_9_2), .weight_en(weight_en));
SA22 U7_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_10_1), .partial_sum_in12(reg_psum6_10_2), .weight_in11(reg_weight6_10_1), .weight_in12(reg_weight6_10_2), .activation_in11(reg_activation7_9_1), .activation_in21(reg_activation7_9_2), .reg_partial_sum21(reg_psum7_10_1), .reg_partial_sum22(reg_psum7_10_2), .reg_weight21(reg_weight7_10_1), .reg_weight22(reg_weight7_10_2), .reg_activation12(reg_activation7_10_1), .reg_activation22(reg_activation7_10_2), .weight_en(weight_en));
SA22 U7_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_11_1), .partial_sum_in12(reg_psum6_11_2), .weight_in11(reg_weight6_11_1), .weight_in12(reg_weight6_11_2), .activation_in11(reg_activation7_10_1), .activation_in21(reg_activation7_10_2), .reg_partial_sum21(reg_psum7_11_1), .reg_partial_sum22(reg_psum7_11_2), .reg_weight21(reg_weight7_11_1), .reg_weight22(reg_weight7_11_2), .reg_activation12(reg_activation7_11_1), .reg_activation22(reg_activation7_11_2), .weight_en(weight_en));
SA22 U7_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_12_1), .partial_sum_in12(reg_psum6_12_2), .weight_in11(reg_weight6_12_1), .weight_in12(reg_weight6_12_2), .activation_in11(reg_activation7_11_1), .activation_in21(reg_activation7_11_2), .reg_partial_sum21(reg_psum7_12_1), .reg_partial_sum22(reg_psum7_12_2), .reg_weight21(reg_weight7_12_1), .reg_weight22(reg_weight7_12_2), .reg_activation12(reg_activation7_12_1), .reg_activation22(reg_activation7_12_2), .weight_en(weight_en));
SA22 U7_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_13_1), .partial_sum_in12(reg_psum6_13_2), .weight_in11(reg_weight6_13_1), .weight_in12(reg_weight6_13_2), .activation_in11(reg_activation7_12_1), .activation_in21(reg_activation7_12_2), .reg_partial_sum21(reg_psum7_13_1), .reg_partial_sum22(reg_psum7_13_2), .reg_weight21(reg_weight7_13_1), .reg_weight22(reg_weight7_13_2), .reg_activation12(reg_activation7_13_1), .reg_activation22(reg_activation7_13_2), .weight_en(weight_en));
SA22 U7_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_14_1), .partial_sum_in12(reg_psum6_14_2), .weight_in11(reg_weight6_14_1), .weight_in12(reg_weight6_14_2), .activation_in11(reg_activation7_13_1), .activation_in21(reg_activation7_13_2), .reg_partial_sum21(reg_psum7_14_1), .reg_partial_sum22(reg_psum7_14_2), .reg_weight21(reg_weight7_14_1), .reg_weight22(reg_weight7_14_2), .reg_activation12(reg_activation7_14_1), .reg_activation22(reg_activation7_14_2), .weight_en(weight_en));
SA22 U7_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_15_1), .partial_sum_in12(reg_psum6_15_2), .weight_in11(reg_weight6_15_1), .weight_in12(reg_weight6_15_2), .activation_in11(reg_activation7_14_1), .activation_in21(reg_activation7_14_2), .reg_partial_sum21(reg_psum7_15_1), .reg_partial_sum22(reg_psum7_15_2), .reg_weight21(reg_weight7_15_1), .reg_weight22(reg_weight7_15_2), .reg_activation12(reg_activation7_15_1), .reg_activation22(reg_activation7_15_2), .weight_en(weight_en));
SA22 U7_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_16_1), .partial_sum_in12(reg_psum6_16_2), .weight_in11(reg_weight6_16_1), .weight_in12(reg_weight6_16_2), .activation_in11(reg_activation7_15_1), .activation_in21(reg_activation7_15_2), .reg_partial_sum21(reg_psum7_16_1), .reg_partial_sum22(reg_psum7_16_2), .reg_weight21(reg_weight7_16_1), .reg_weight22(reg_weight7_16_2), .reg_activation12(reg_activation7_16_1), .reg_activation22(reg_activation7_16_2), .weight_en(weight_en));
SA22 U7_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_17_1), .partial_sum_in12(reg_psum6_17_2), .weight_in11(reg_weight6_17_1), .weight_in12(reg_weight6_17_2), .activation_in11(reg_activation7_16_1), .activation_in21(reg_activation7_16_2), .reg_partial_sum21(reg_psum7_17_1), .reg_partial_sum22(reg_psum7_17_2), .reg_weight21(reg_weight7_17_1), .reg_weight22(reg_weight7_17_2), .reg_activation12(reg_activation7_17_1), .reg_activation22(reg_activation7_17_2), .weight_en(weight_en));
SA22 U7_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_18_1), .partial_sum_in12(reg_psum6_18_2), .weight_in11(reg_weight6_18_1), .weight_in12(reg_weight6_18_2), .activation_in11(reg_activation7_17_1), .activation_in21(reg_activation7_17_2), .reg_partial_sum21(reg_psum7_18_1), .reg_partial_sum22(reg_psum7_18_2), .reg_weight21(reg_weight7_18_1), .reg_weight22(reg_weight7_18_2), .reg_activation12(reg_activation7_18_1), .reg_activation22(reg_activation7_18_2), .weight_en(weight_en));
SA22 U7_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_19_1), .partial_sum_in12(reg_psum6_19_2), .weight_in11(reg_weight6_19_1), .weight_in12(reg_weight6_19_2), .activation_in11(reg_activation7_18_1), .activation_in21(reg_activation7_18_2), .reg_partial_sum21(reg_psum7_19_1), .reg_partial_sum22(reg_psum7_19_2), .reg_weight21(reg_weight7_19_1), .reg_weight22(reg_weight7_19_2), .reg_activation12(reg_activation7_19_1), .reg_activation22(reg_activation7_19_2), .weight_en(weight_en));
SA22 U7_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_20_1), .partial_sum_in12(reg_psum6_20_2), .weight_in11(reg_weight6_20_1), .weight_in12(reg_weight6_20_2), .activation_in11(reg_activation7_19_1), .activation_in21(reg_activation7_19_2), .reg_partial_sum21(reg_psum7_20_1), .reg_partial_sum22(reg_psum7_20_2), .reg_weight21(reg_weight7_20_1), .reg_weight22(reg_weight7_20_2), .reg_activation12(reg_activation7_20_1), .reg_activation22(reg_activation7_20_2), .weight_en(weight_en));
SA22 U7_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_21_1), .partial_sum_in12(reg_psum6_21_2), .weight_in11(reg_weight6_21_1), .weight_in12(reg_weight6_21_2), .activation_in11(reg_activation7_20_1), .activation_in21(reg_activation7_20_2), .reg_partial_sum21(reg_psum7_21_1), .reg_partial_sum22(reg_psum7_21_2), .reg_weight21(reg_weight7_21_1), .reg_weight22(reg_weight7_21_2), .reg_activation12(reg_activation7_21_1), .reg_activation22(reg_activation7_21_2), .weight_en(weight_en));
SA22 U7_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_22_1), .partial_sum_in12(reg_psum6_22_2), .weight_in11(reg_weight6_22_1), .weight_in12(reg_weight6_22_2), .activation_in11(reg_activation7_21_1), .activation_in21(reg_activation7_21_2), .reg_partial_sum21(reg_psum7_22_1), .reg_partial_sum22(reg_psum7_22_2), .reg_weight21(reg_weight7_22_1), .reg_weight22(reg_weight7_22_2), .reg_activation12(reg_activation7_22_1), .reg_activation22(reg_activation7_22_2), .weight_en(weight_en));
SA22 U7_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_23_1), .partial_sum_in12(reg_psum6_23_2), .weight_in11(reg_weight6_23_1), .weight_in12(reg_weight6_23_2), .activation_in11(reg_activation7_22_1), .activation_in21(reg_activation7_22_2), .reg_partial_sum21(reg_psum7_23_1), .reg_partial_sum22(reg_psum7_23_2), .reg_weight21(reg_weight7_23_1), .reg_weight22(reg_weight7_23_2), .reg_activation12(reg_activation7_23_1), .reg_activation22(reg_activation7_23_2), .weight_en(weight_en));
SA22 U7_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_24_1), .partial_sum_in12(reg_psum6_24_2), .weight_in11(reg_weight6_24_1), .weight_in12(reg_weight6_24_2), .activation_in11(reg_activation7_23_1), .activation_in21(reg_activation7_23_2), .reg_partial_sum21(reg_psum7_24_1), .reg_partial_sum22(reg_psum7_24_2), .reg_weight21(reg_weight7_24_1), .reg_weight22(reg_weight7_24_2), .reg_activation12(reg_activation7_24_1), .reg_activation22(reg_activation7_24_2), .weight_en(weight_en));
SA22 U7_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_25_1), .partial_sum_in12(reg_psum6_25_2), .weight_in11(reg_weight6_25_1), .weight_in12(reg_weight6_25_2), .activation_in11(reg_activation7_24_1), .activation_in21(reg_activation7_24_2), .reg_partial_sum21(reg_psum7_25_1), .reg_partial_sum22(reg_psum7_25_2), .reg_weight21(reg_weight7_25_1), .reg_weight22(reg_weight7_25_2), .reg_activation12(reg_activation7_25_1), .reg_activation22(reg_activation7_25_2), .weight_en(weight_en));
SA22 U7_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_26_1), .partial_sum_in12(reg_psum6_26_2), .weight_in11(reg_weight6_26_1), .weight_in12(reg_weight6_26_2), .activation_in11(reg_activation7_25_1), .activation_in21(reg_activation7_25_2), .reg_partial_sum21(reg_psum7_26_1), .reg_partial_sum22(reg_psum7_26_2), .reg_weight21(reg_weight7_26_1), .reg_weight22(reg_weight7_26_2), .reg_activation12(reg_activation7_26_1), .reg_activation22(reg_activation7_26_2), .weight_en(weight_en));
SA22 U7_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_27_1), .partial_sum_in12(reg_psum6_27_2), .weight_in11(reg_weight6_27_1), .weight_in12(reg_weight6_27_2), .activation_in11(reg_activation7_26_1), .activation_in21(reg_activation7_26_2), .reg_partial_sum21(reg_psum7_27_1), .reg_partial_sum22(reg_psum7_27_2), .reg_weight21(reg_weight7_27_1), .reg_weight22(reg_weight7_27_2), .reg_activation12(reg_activation7_27_1), .reg_activation22(reg_activation7_27_2), .weight_en(weight_en));
SA22 U7_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_28_1), .partial_sum_in12(reg_psum6_28_2), .weight_in11(reg_weight6_28_1), .weight_in12(reg_weight6_28_2), .activation_in11(reg_activation7_27_1), .activation_in21(reg_activation7_27_2), .reg_partial_sum21(reg_psum7_28_1), .reg_partial_sum22(reg_psum7_28_2), .reg_weight21(reg_weight7_28_1), .reg_weight22(reg_weight7_28_2), .reg_activation12(reg_activation7_28_1), .reg_activation22(reg_activation7_28_2), .weight_en(weight_en));
SA22 U7_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_29_1), .partial_sum_in12(reg_psum6_29_2), .weight_in11(reg_weight6_29_1), .weight_in12(reg_weight6_29_2), .activation_in11(reg_activation7_28_1), .activation_in21(reg_activation7_28_2), .reg_partial_sum21(reg_psum7_29_1), .reg_partial_sum22(reg_psum7_29_2), .reg_weight21(reg_weight7_29_1), .reg_weight22(reg_weight7_29_2), .reg_activation12(reg_activation7_29_1), .reg_activation22(reg_activation7_29_2), .weight_en(weight_en));
SA22 U7_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_30_1), .partial_sum_in12(reg_psum6_30_2), .weight_in11(reg_weight6_30_1), .weight_in12(reg_weight6_30_2), .activation_in11(reg_activation7_29_1), .activation_in21(reg_activation7_29_2), .reg_partial_sum21(reg_psum7_30_1), .reg_partial_sum22(reg_psum7_30_2), .reg_weight21(reg_weight7_30_1), .reg_weight22(reg_weight7_30_2), .reg_activation12(reg_activation7_30_1), .reg_activation22(reg_activation7_30_2), .weight_en(weight_en));
SA22 U7_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_31_1), .partial_sum_in12(reg_psum6_31_2), .weight_in11(reg_weight6_31_1), .weight_in12(reg_weight6_31_2), .activation_in11(reg_activation7_30_1), .activation_in21(reg_activation7_30_2), .reg_partial_sum21(reg_psum7_31_1), .reg_partial_sum22(reg_psum7_31_2), .reg_weight21(reg_weight7_31_1), .reg_weight22(reg_weight7_31_2), .reg_activation12(reg_activation7_31_1), .reg_activation22(reg_activation7_31_2), .weight_en(weight_en));
SA22 U7_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum6_32_1), .partial_sum_in12(reg_psum6_32_2), .weight_in11(reg_weight6_32_1), .weight_in12(reg_weight6_32_2), .activation_in11(reg_activation7_31_1), .activation_in21(reg_activation7_31_2), .reg_partial_sum21(reg_psum7_32_1), .reg_partial_sum22(reg_psum7_32_2), .reg_weight21(reg_weight7_32_1), .reg_weight22(reg_weight7_32_2), .weight_en(weight_en));
SA22 U8_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_1_1), .partial_sum_in12(reg_psum7_1_2), .weight_in11(reg_weight7_1_1), .weight_in12(reg_weight7_1_2), .activation_in11(in_activation8_1_1), .activation_in21(in_activation8_1_2), .reg_partial_sum21(reg_psum8_1_1), .reg_partial_sum22(reg_psum8_1_2), .reg_weight21(reg_weight8_1_1), .reg_weight22(reg_weight8_1_2), .reg_activation12(reg_activation8_1_1), .reg_activation22(reg_activation8_1_2), .weight_en(weight_en));
SA22 U8_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_2_1), .partial_sum_in12(reg_psum7_2_2), .weight_in11(reg_weight7_2_1), .weight_in12(reg_weight7_2_2), .activation_in11(reg_activation8_1_1), .activation_in21(reg_activation8_1_2), .reg_partial_sum21(reg_psum8_2_1), .reg_partial_sum22(reg_psum8_2_2), .reg_weight21(reg_weight8_2_1), .reg_weight22(reg_weight8_2_2), .reg_activation12(reg_activation8_2_1), .reg_activation22(reg_activation8_2_2), .weight_en(weight_en));
SA22 U8_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_3_1), .partial_sum_in12(reg_psum7_3_2), .weight_in11(reg_weight7_3_1), .weight_in12(reg_weight7_3_2), .activation_in11(reg_activation8_2_1), .activation_in21(reg_activation8_2_2), .reg_partial_sum21(reg_psum8_3_1), .reg_partial_sum22(reg_psum8_3_2), .reg_weight21(reg_weight8_3_1), .reg_weight22(reg_weight8_3_2), .reg_activation12(reg_activation8_3_1), .reg_activation22(reg_activation8_3_2), .weight_en(weight_en));
SA22 U8_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_4_1), .partial_sum_in12(reg_psum7_4_2), .weight_in11(reg_weight7_4_1), .weight_in12(reg_weight7_4_2), .activation_in11(reg_activation8_3_1), .activation_in21(reg_activation8_3_2), .reg_partial_sum21(reg_psum8_4_1), .reg_partial_sum22(reg_psum8_4_2), .reg_weight21(reg_weight8_4_1), .reg_weight22(reg_weight8_4_2), .reg_activation12(reg_activation8_4_1), .reg_activation22(reg_activation8_4_2), .weight_en(weight_en));
SA22 U8_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_5_1), .partial_sum_in12(reg_psum7_5_2), .weight_in11(reg_weight7_5_1), .weight_in12(reg_weight7_5_2), .activation_in11(reg_activation8_4_1), .activation_in21(reg_activation8_4_2), .reg_partial_sum21(reg_psum8_5_1), .reg_partial_sum22(reg_psum8_5_2), .reg_weight21(reg_weight8_5_1), .reg_weight22(reg_weight8_5_2), .reg_activation12(reg_activation8_5_1), .reg_activation22(reg_activation8_5_2), .weight_en(weight_en));
SA22 U8_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_6_1), .partial_sum_in12(reg_psum7_6_2), .weight_in11(reg_weight7_6_1), .weight_in12(reg_weight7_6_2), .activation_in11(reg_activation8_5_1), .activation_in21(reg_activation8_5_2), .reg_partial_sum21(reg_psum8_6_1), .reg_partial_sum22(reg_psum8_6_2), .reg_weight21(reg_weight8_6_1), .reg_weight22(reg_weight8_6_2), .reg_activation12(reg_activation8_6_1), .reg_activation22(reg_activation8_6_2), .weight_en(weight_en));
SA22 U8_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_7_1), .partial_sum_in12(reg_psum7_7_2), .weight_in11(reg_weight7_7_1), .weight_in12(reg_weight7_7_2), .activation_in11(reg_activation8_6_1), .activation_in21(reg_activation8_6_2), .reg_partial_sum21(reg_psum8_7_1), .reg_partial_sum22(reg_psum8_7_2), .reg_weight21(reg_weight8_7_1), .reg_weight22(reg_weight8_7_2), .reg_activation12(reg_activation8_7_1), .reg_activation22(reg_activation8_7_2), .weight_en(weight_en));
SA22 U8_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_8_1), .partial_sum_in12(reg_psum7_8_2), .weight_in11(reg_weight7_8_1), .weight_in12(reg_weight7_8_2), .activation_in11(reg_activation8_7_1), .activation_in21(reg_activation8_7_2), .reg_partial_sum21(reg_psum8_8_1), .reg_partial_sum22(reg_psum8_8_2), .reg_weight21(reg_weight8_8_1), .reg_weight22(reg_weight8_8_2), .reg_activation12(reg_activation8_8_1), .reg_activation22(reg_activation8_8_2), .weight_en(weight_en));
SA22 U8_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_9_1), .partial_sum_in12(reg_psum7_9_2), .weight_in11(reg_weight7_9_1), .weight_in12(reg_weight7_9_2), .activation_in11(reg_activation8_8_1), .activation_in21(reg_activation8_8_2), .reg_partial_sum21(reg_psum8_9_1), .reg_partial_sum22(reg_psum8_9_2), .reg_weight21(reg_weight8_9_1), .reg_weight22(reg_weight8_9_2), .reg_activation12(reg_activation8_9_1), .reg_activation22(reg_activation8_9_2), .weight_en(weight_en));
SA22 U8_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_10_1), .partial_sum_in12(reg_psum7_10_2), .weight_in11(reg_weight7_10_1), .weight_in12(reg_weight7_10_2), .activation_in11(reg_activation8_9_1), .activation_in21(reg_activation8_9_2), .reg_partial_sum21(reg_psum8_10_1), .reg_partial_sum22(reg_psum8_10_2), .reg_weight21(reg_weight8_10_1), .reg_weight22(reg_weight8_10_2), .reg_activation12(reg_activation8_10_1), .reg_activation22(reg_activation8_10_2), .weight_en(weight_en));
SA22 U8_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_11_1), .partial_sum_in12(reg_psum7_11_2), .weight_in11(reg_weight7_11_1), .weight_in12(reg_weight7_11_2), .activation_in11(reg_activation8_10_1), .activation_in21(reg_activation8_10_2), .reg_partial_sum21(reg_psum8_11_1), .reg_partial_sum22(reg_psum8_11_2), .reg_weight21(reg_weight8_11_1), .reg_weight22(reg_weight8_11_2), .reg_activation12(reg_activation8_11_1), .reg_activation22(reg_activation8_11_2), .weight_en(weight_en));
SA22 U8_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_12_1), .partial_sum_in12(reg_psum7_12_2), .weight_in11(reg_weight7_12_1), .weight_in12(reg_weight7_12_2), .activation_in11(reg_activation8_11_1), .activation_in21(reg_activation8_11_2), .reg_partial_sum21(reg_psum8_12_1), .reg_partial_sum22(reg_psum8_12_2), .reg_weight21(reg_weight8_12_1), .reg_weight22(reg_weight8_12_2), .reg_activation12(reg_activation8_12_1), .reg_activation22(reg_activation8_12_2), .weight_en(weight_en));
SA22 U8_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_13_1), .partial_sum_in12(reg_psum7_13_2), .weight_in11(reg_weight7_13_1), .weight_in12(reg_weight7_13_2), .activation_in11(reg_activation8_12_1), .activation_in21(reg_activation8_12_2), .reg_partial_sum21(reg_psum8_13_1), .reg_partial_sum22(reg_psum8_13_2), .reg_weight21(reg_weight8_13_1), .reg_weight22(reg_weight8_13_2), .reg_activation12(reg_activation8_13_1), .reg_activation22(reg_activation8_13_2), .weight_en(weight_en));
SA22 U8_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_14_1), .partial_sum_in12(reg_psum7_14_2), .weight_in11(reg_weight7_14_1), .weight_in12(reg_weight7_14_2), .activation_in11(reg_activation8_13_1), .activation_in21(reg_activation8_13_2), .reg_partial_sum21(reg_psum8_14_1), .reg_partial_sum22(reg_psum8_14_2), .reg_weight21(reg_weight8_14_1), .reg_weight22(reg_weight8_14_2), .reg_activation12(reg_activation8_14_1), .reg_activation22(reg_activation8_14_2), .weight_en(weight_en));
SA22 U8_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_15_1), .partial_sum_in12(reg_psum7_15_2), .weight_in11(reg_weight7_15_1), .weight_in12(reg_weight7_15_2), .activation_in11(reg_activation8_14_1), .activation_in21(reg_activation8_14_2), .reg_partial_sum21(reg_psum8_15_1), .reg_partial_sum22(reg_psum8_15_2), .reg_weight21(reg_weight8_15_1), .reg_weight22(reg_weight8_15_2), .reg_activation12(reg_activation8_15_1), .reg_activation22(reg_activation8_15_2), .weight_en(weight_en));
SA22 U8_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_16_1), .partial_sum_in12(reg_psum7_16_2), .weight_in11(reg_weight7_16_1), .weight_in12(reg_weight7_16_2), .activation_in11(reg_activation8_15_1), .activation_in21(reg_activation8_15_2), .reg_partial_sum21(reg_psum8_16_1), .reg_partial_sum22(reg_psum8_16_2), .reg_weight21(reg_weight8_16_1), .reg_weight22(reg_weight8_16_2), .reg_activation12(reg_activation8_16_1), .reg_activation22(reg_activation8_16_2), .weight_en(weight_en));
SA22 U8_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_17_1), .partial_sum_in12(reg_psum7_17_2), .weight_in11(reg_weight7_17_1), .weight_in12(reg_weight7_17_2), .activation_in11(reg_activation8_16_1), .activation_in21(reg_activation8_16_2), .reg_partial_sum21(reg_psum8_17_1), .reg_partial_sum22(reg_psum8_17_2), .reg_weight21(reg_weight8_17_1), .reg_weight22(reg_weight8_17_2), .reg_activation12(reg_activation8_17_1), .reg_activation22(reg_activation8_17_2), .weight_en(weight_en));
SA22 U8_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_18_1), .partial_sum_in12(reg_psum7_18_2), .weight_in11(reg_weight7_18_1), .weight_in12(reg_weight7_18_2), .activation_in11(reg_activation8_17_1), .activation_in21(reg_activation8_17_2), .reg_partial_sum21(reg_psum8_18_1), .reg_partial_sum22(reg_psum8_18_2), .reg_weight21(reg_weight8_18_1), .reg_weight22(reg_weight8_18_2), .reg_activation12(reg_activation8_18_1), .reg_activation22(reg_activation8_18_2), .weight_en(weight_en));
SA22 U8_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_19_1), .partial_sum_in12(reg_psum7_19_2), .weight_in11(reg_weight7_19_1), .weight_in12(reg_weight7_19_2), .activation_in11(reg_activation8_18_1), .activation_in21(reg_activation8_18_2), .reg_partial_sum21(reg_psum8_19_1), .reg_partial_sum22(reg_psum8_19_2), .reg_weight21(reg_weight8_19_1), .reg_weight22(reg_weight8_19_2), .reg_activation12(reg_activation8_19_1), .reg_activation22(reg_activation8_19_2), .weight_en(weight_en));
SA22 U8_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_20_1), .partial_sum_in12(reg_psum7_20_2), .weight_in11(reg_weight7_20_1), .weight_in12(reg_weight7_20_2), .activation_in11(reg_activation8_19_1), .activation_in21(reg_activation8_19_2), .reg_partial_sum21(reg_psum8_20_1), .reg_partial_sum22(reg_psum8_20_2), .reg_weight21(reg_weight8_20_1), .reg_weight22(reg_weight8_20_2), .reg_activation12(reg_activation8_20_1), .reg_activation22(reg_activation8_20_2), .weight_en(weight_en));
SA22 U8_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_21_1), .partial_sum_in12(reg_psum7_21_2), .weight_in11(reg_weight7_21_1), .weight_in12(reg_weight7_21_2), .activation_in11(reg_activation8_20_1), .activation_in21(reg_activation8_20_2), .reg_partial_sum21(reg_psum8_21_1), .reg_partial_sum22(reg_psum8_21_2), .reg_weight21(reg_weight8_21_1), .reg_weight22(reg_weight8_21_2), .reg_activation12(reg_activation8_21_1), .reg_activation22(reg_activation8_21_2), .weight_en(weight_en));
SA22 U8_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_22_1), .partial_sum_in12(reg_psum7_22_2), .weight_in11(reg_weight7_22_1), .weight_in12(reg_weight7_22_2), .activation_in11(reg_activation8_21_1), .activation_in21(reg_activation8_21_2), .reg_partial_sum21(reg_psum8_22_1), .reg_partial_sum22(reg_psum8_22_2), .reg_weight21(reg_weight8_22_1), .reg_weight22(reg_weight8_22_2), .reg_activation12(reg_activation8_22_1), .reg_activation22(reg_activation8_22_2), .weight_en(weight_en));
SA22 U8_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_23_1), .partial_sum_in12(reg_psum7_23_2), .weight_in11(reg_weight7_23_1), .weight_in12(reg_weight7_23_2), .activation_in11(reg_activation8_22_1), .activation_in21(reg_activation8_22_2), .reg_partial_sum21(reg_psum8_23_1), .reg_partial_sum22(reg_psum8_23_2), .reg_weight21(reg_weight8_23_1), .reg_weight22(reg_weight8_23_2), .reg_activation12(reg_activation8_23_1), .reg_activation22(reg_activation8_23_2), .weight_en(weight_en));
SA22 U8_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_24_1), .partial_sum_in12(reg_psum7_24_2), .weight_in11(reg_weight7_24_1), .weight_in12(reg_weight7_24_2), .activation_in11(reg_activation8_23_1), .activation_in21(reg_activation8_23_2), .reg_partial_sum21(reg_psum8_24_1), .reg_partial_sum22(reg_psum8_24_2), .reg_weight21(reg_weight8_24_1), .reg_weight22(reg_weight8_24_2), .reg_activation12(reg_activation8_24_1), .reg_activation22(reg_activation8_24_2), .weight_en(weight_en));
SA22 U8_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_25_1), .partial_sum_in12(reg_psum7_25_2), .weight_in11(reg_weight7_25_1), .weight_in12(reg_weight7_25_2), .activation_in11(reg_activation8_24_1), .activation_in21(reg_activation8_24_2), .reg_partial_sum21(reg_psum8_25_1), .reg_partial_sum22(reg_psum8_25_2), .reg_weight21(reg_weight8_25_1), .reg_weight22(reg_weight8_25_2), .reg_activation12(reg_activation8_25_1), .reg_activation22(reg_activation8_25_2), .weight_en(weight_en));
SA22 U8_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_26_1), .partial_sum_in12(reg_psum7_26_2), .weight_in11(reg_weight7_26_1), .weight_in12(reg_weight7_26_2), .activation_in11(reg_activation8_25_1), .activation_in21(reg_activation8_25_2), .reg_partial_sum21(reg_psum8_26_1), .reg_partial_sum22(reg_psum8_26_2), .reg_weight21(reg_weight8_26_1), .reg_weight22(reg_weight8_26_2), .reg_activation12(reg_activation8_26_1), .reg_activation22(reg_activation8_26_2), .weight_en(weight_en));
SA22 U8_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_27_1), .partial_sum_in12(reg_psum7_27_2), .weight_in11(reg_weight7_27_1), .weight_in12(reg_weight7_27_2), .activation_in11(reg_activation8_26_1), .activation_in21(reg_activation8_26_2), .reg_partial_sum21(reg_psum8_27_1), .reg_partial_sum22(reg_psum8_27_2), .reg_weight21(reg_weight8_27_1), .reg_weight22(reg_weight8_27_2), .reg_activation12(reg_activation8_27_1), .reg_activation22(reg_activation8_27_2), .weight_en(weight_en));
SA22 U8_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_28_1), .partial_sum_in12(reg_psum7_28_2), .weight_in11(reg_weight7_28_1), .weight_in12(reg_weight7_28_2), .activation_in11(reg_activation8_27_1), .activation_in21(reg_activation8_27_2), .reg_partial_sum21(reg_psum8_28_1), .reg_partial_sum22(reg_psum8_28_2), .reg_weight21(reg_weight8_28_1), .reg_weight22(reg_weight8_28_2), .reg_activation12(reg_activation8_28_1), .reg_activation22(reg_activation8_28_2), .weight_en(weight_en));
SA22 U8_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_29_1), .partial_sum_in12(reg_psum7_29_2), .weight_in11(reg_weight7_29_1), .weight_in12(reg_weight7_29_2), .activation_in11(reg_activation8_28_1), .activation_in21(reg_activation8_28_2), .reg_partial_sum21(reg_psum8_29_1), .reg_partial_sum22(reg_psum8_29_2), .reg_weight21(reg_weight8_29_1), .reg_weight22(reg_weight8_29_2), .reg_activation12(reg_activation8_29_1), .reg_activation22(reg_activation8_29_2), .weight_en(weight_en));
SA22 U8_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_30_1), .partial_sum_in12(reg_psum7_30_2), .weight_in11(reg_weight7_30_1), .weight_in12(reg_weight7_30_2), .activation_in11(reg_activation8_29_1), .activation_in21(reg_activation8_29_2), .reg_partial_sum21(reg_psum8_30_1), .reg_partial_sum22(reg_psum8_30_2), .reg_weight21(reg_weight8_30_1), .reg_weight22(reg_weight8_30_2), .reg_activation12(reg_activation8_30_1), .reg_activation22(reg_activation8_30_2), .weight_en(weight_en));
SA22 U8_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_31_1), .partial_sum_in12(reg_psum7_31_2), .weight_in11(reg_weight7_31_1), .weight_in12(reg_weight7_31_2), .activation_in11(reg_activation8_30_1), .activation_in21(reg_activation8_30_2), .reg_partial_sum21(reg_psum8_31_1), .reg_partial_sum22(reg_psum8_31_2), .reg_weight21(reg_weight8_31_1), .reg_weight22(reg_weight8_31_2), .reg_activation12(reg_activation8_31_1), .reg_activation22(reg_activation8_31_2), .weight_en(weight_en));
SA22 U8_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum7_32_1), .partial_sum_in12(reg_psum7_32_2), .weight_in11(reg_weight7_32_1), .weight_in12(reg_weight7_32_2), .activation_in11(reg_activation8_31_1), .activation_in21(reg_activation8_31_2), .reg_partial_sum21(reg_psum8_32_1), .reg_partial_sum22(reg_psum8_32_2), .reg_weight21(reg_weight8_32_1), .reg_weight22(reg_weight8_32_2), .weight_en(weight_en));
SA22 U9_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_1_1), .partial_sum_in12(reg_psum8_1_2), .weight_in11(reg_weight8_1_1), .weight_in12(reg_weight8_1_2), .activation_in11(in_activation9_1_1), .activation_in21(in_activation9_1_2), .reg_partial_sum21(reg_psum9_1_1), .reg_partial_sum22(reg_psum9_1_2), .reg_weight21(reg_weight9_1_1), .reg_weight22(reg_weight9_1_2), .reg_activation12(reg_activation9_1_1), .reg_activation22(reg_activation9_1_2), .weight_en(weight_en));
SA22 U9_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_2_1), .partial_sum_in12(reg_psum8_2_2), .weight_in11(reg_weight8_2_1), .weight_in12(reg_weight8_2_2), .activation_in11(reg_activation9_1_1), .activation_in21(reg_activation9_1_2), .reg_partial_sum21(reg_psum9_2_1), .reg_partial_sum22(reg_psum9_2_2), .reg_weight21(reg_weight9_2_1), .reg_weight22(reg_weight9_2_2), .reg_activation12(reg_activation9_2_1), .reg_activation22(reg_activation9_2_2), .weight_en(weight_en));
SA22 U9_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_3_1), .partial_sum_in12(reg_psum8_3_2), .weight_in11(reg_weight8_3_1), .weight_in12(reg_weight8_3_2), .activation_in11(reg_activation9_2_1), .activation_in21(reg_activation9_2_2), .reg_partial_sum21(reg_psum9_3_1), .reg_partial_sum22(reg_psum9_3_2), .reg_weight21(reg_weight9_3_1), .reg_weight22(reg_weight9_3_2), .reg_activation12(reg_activation9_3_1), .reg_activation22(reg_activation9_3_2), .weight_en(weight_en));
SA22 U9_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_4_1), .partial_sum_in12(reg_psum8_4_2), .weight_in11(reg_weight8_4_1), .weight_in12(reg_weight8_4_2), .activation_in11(reg_activation9_3_1), .activation_in21(reg_activation9_3_2), .reg_partial_sum21(reg_psum9_4_1), .reg_partial_sum22(reg_psum9_4_2), .reg_weight21(reg_weight9_4_1), .reg_weight22(reg_weight9_4_2), .reg_activation12(reg_activation9_4_1), .reg_activation22(reg_activation9_4_2), .weight_en(weight_en));
SA22 U9_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_5_1), .partial_sum_in12(reg_psum8_5_2), .weight_in11(reg_weight8_5_1), .weight_in12(reg_weight8_5_2), .activation_in11(reg_activation9_4_1), .activation_in21(reg_activation9_4_2), .reg_partial_sum21(reg_psum9_5_1), .reg_partial_sum22(reg_psum9_5_2), .reg_weight21(reg_weight9_5_1), .reg_weight22(reg_weight9_5_2), .reg_activation12(reg_activation9_5_1), .reg_activation22(reg_activation9_5_2), .weight_en(weight_en));
SA22 U9_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_6_1), .partial_sum_in12(reg_psum8_6_2), .weight_in11(reg_weight8_6_1), .weight_in12(reg_weight8_6_2), .activation_in11(reg_activation9_5_1), .activation_in21(reg_activation9_5_2), .reg_partial_sum21(reg_psum9_6_1), .reg_partial_sum22(reg_psum9_6_2), .reg_weight21(reg_weight9_6_1), .reg_weight22(reg_weight9_6_2), .reg_activation12(reg_activation9_6_1), .reg_activation22(reg_activation9_6_2), .weight_en(weight_en));
SA22 U9_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_7_1), .partial_sum_in12(reg_psum8_7_2), .weight_in11(reg_weight8_7_1), .weight_in12(reg_weight8_7_2), .activation_in11(reg_activation9_6_1), .activation_in21(reg_activation9_6_2), .reg_partial_sum21(reg_psum9_7_1), .reg_partial_sum22(reg_psum9_7_2), .reg_weight21(reg_weight9_7_1), .reg_weight22(reg_weight9_7_2), .reg_activation12(reg_activation9_7_1), .reg_activation22(reg_activation9_7_2), .weight_en(weight_en));
SA22 U9_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_8_1), .partial_sum_in12(reg_psum8_8_2), .weight_in11(reg_weight8_8_1), .weight_in12(reg_weight8_8_2), .activation_in11(reg_activation9_7_1), .activation_in21(reg_activation9_7_2), .reg_partial_sum21(reg_psum9_8_1), .reg_partial_sum22(reg_psum9_8_2), .reg_weight21(reg_weight9_8_1), .reg_weight22(reg_weight9_8_2), .reg_activation12(reg_activation9_8_1), .reg_activation22(reg_activation9_8_2), .weight_en(weight_en));
SA22 U9_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_9_1), .partial_sum_in12(reg_psum8_9_2), .weight_in11(reg_weight8_9_1), .weight_in12(reg_weight8_9_2), .activation_in11(reg_activation9_8_1), .activation_in21(reg_activation9_8_2), .reg_partial_sum21(reg_psum9_9_1), .reg_partial_sum22(reg_psum9_9_2), .reg_weight21(reg_weight9_9_1), .reg_weight22(reg_weight9_9_2), .reg_activation12(reg_activation9_9_1), .reg_activation22(reg_activation9_9_2), .weight_en(weight_en));
SA22 U9_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_10_1), .partial_sum_in12(reg_psum8_10_2), .weight_in11(reg_weight8_10_1), .weight_in12(reg_weight8_10_2), .activation_in11(reg_activation9_9_1), .activation_in21(reg_activation9_9_2), .reg_partial_sum21(reg_psum9_10_1), .reg_partial_sum22(reg_psum9_10_2), .reg_weight21(reg_weight9_10_1), .reg_weight22(reg_weight9_10_2), .reg_activation12(reg_activation9_10_1), .reg_activation22(reg_activation9_10_2), .weight_en(weight_en));
SA22 U9_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_11_1), .partial_sum_in12(reg_psum8_11_2), .weight_in11(reg_weight8_11_1), .weight_in12(reg_weight8_11_2), .activation_in11(reg_activation9_10_1), .activation_in21(reg_activation9_10_2), .reg_partial_sum21(reg_psum9_11_1), .reg_partial_sum22(reg_psum9_11_2), .reg_weight21(reg_weight9_11_1), .reg_weight22(reg_weight9_11_2), .reg_activation12(reg_activation9_11_1), .reg_activation22(reg_activation9_11_2), .weight_en(weight_en));
SA22 U9_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_12_1), .partial_sum_in12(reg_psum8_12_2), .weight_in11(reg_weight8_12_1), .weight_in12(reg_weight8_12_2), .activation_in11(reg_activation9_11_1), .activation_in21(reg_activation9_11_2), .reg_partial_sum21(reg_psum9_12_1), .reg_partial_sum22(reg_psum9_12_2), .reg_weight21(reg_weight9_12_1), .reg_weight22(reg_weight9_12_2), .reg_activation12(reg_activation9_12_1), .reg_activation22(reg_activation9_12_2), .weight_en(weight_en));
SA22 U9_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_13_1), .partial_sum_in12(reg_psum8_13_2), .weight_in11(reg_weight8_13_1), .weight_in12(reg_weight8_13_2), .activation_in11(reg_activation9_12_1), .activation_in21(reg_activation9_12_2), .reg_partial_sum21(reg_psum9_13_1), .reg_partial_sum22(reg_psum9_13_2), .reg_weight21(reg_weight9_13_1), .reg_weight22(reg_weight9_13_2), .reg_activation12(reg_activation9_13_1), .reg_activation22(reg_activation9_13_2), .weight_en(weight_en));
SA22 U9_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_14_1), .partial_sum_in12(reg_psum8_14_2), .weight_in11(reg_weight8_14_1), .weight_in12(reg_weight8_14_2), .activation_in11(reg_activation9_13_1), .activation_in21(reg_activation9_13_2), .reg_partial_sum21(reg_psum9_14_1), .reg_partial_sum22(reg_psum9_14_2), .reg_weight21(reg_weight9_14_1), .reg_weight22(reg_weight9_14_2), .reg_activation12(reg_activation9_14_1), .reg_activation22(reg_activation9_14_2), .weight_en(weight_en));
SA22 U9_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_15_1), .partial_sum_in12(reg_psum8_15_2), .weight_in11(reg_weight8_15_1), .weight_in12(reg_weight8_15_2), .activation_in11(reg_activation9_14_1), .activation_in21(reg_activation9_14_2), .reg_partial_sum21(reg_psum9_15_1), .reg_partial_sum22(reg_psum9_15_2), .reg_weight21(reg_weight9_15_1), .reg_weight22(reg_weight9_15_2), .reg_activation12(reg_activation9_15_1), .reg_activation22(reg_activation9_15_2), .weight_en(weight_en));
SA22 U9_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_16_1), .partial_sum_in12(reg_psum8_16_2), .weight_in11(reg_weight8_16_1), .weight_in12(reg_weight8_16_2), .activation_in11(reg_activation9_15_1), .activation_in21(reg_activation9_15_2), .reg_partial_sum21(reg_psum9_16_1), .reg_partial_sum22(reg_psum9_16_2), .reg_weight21(reg_weight9_16_1), .reg_weight22(reg_weight9_16_2), .reg_activation12(reg_activation9_16_1), .reg_activation22(reg_activation9_16_2), .weight_en(weight_en));
SA22 U9_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_17_1), .partial_sum_in12(reg_psum8_17_2), .weight_in11(reg_weight8_17_1), .weight_in12(reg_weight8_17_2), .activation_in11(reg_activation9_16_1), .activation_in21(reg_activation9_16_2), .reg_partial_sum21(reg_psum9_17_1), .reg_partial_sum22(reg_psum9_17_2), .reg_weight21(reg_weight9_17_1), .reg_weight22(reg_weight9_17_2), .reg_activation12(reg_activation9_17_1), .reg_activation22(reg_activation9_17_2), .weight_en(weight_en));
SA22 U9_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_18_1), .partial_sum_in12(reg_psum8_18_2), .weight_in11(reg_weight8_18_1), .weight_in12(reg_weight8_18_2), .activation_in11(reg_activation9_17_1), .activation_in21(reg_activation9_17_2), .reg_partial_sum21(reg_psum9_18_1), .reg_partial_sum22(reg_psum9_18_2), .reg_weight21(reg_weight9_18_1), .reg_weight22(reg_weight9_18_2), .reg_activation12(reg_activation9_18_1), .reg_activation22(reg_activation9_18_2), .weight_en(weight_en));
SA22 U9_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_19_1), .partial_sum_in12(reg_psum8_19_2), .weight_in11(reg_weight8_19_1), .weight_in12(reg_weight8_19_2), .activation_in11(reg_activation9_18_1), .activation_in21(reg_activation9_18_2), .reg_partial_sum21(reg_psum9_19_1), .reg_partial_sum22(reg_psum9_19_2), .reg_weight21(reg_weight9_19_1), .reg_weight22(reg_weight9_19_2), .reg_activation12(reg_activation9_19_1), .reg_activation22(reg_activation9_19_2), .weight_en(weight_en));
SA22 U9_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_20_1), .partial_sum_in12(reg_psum8_20_2), .weight_in11(reg_weight8_20_1), .weight_in12(reg_weight8_20_2), .activation_in11(reg_activation9_19_1), .activation_in21(reg_activation9_19_2), .reg_partial_sum21(reg_psum9_20_1), .reg_partial_sum22(reg_psum9_20_2), .reg_weight21(reg_weight9_20_1), .reg_weight22(reg_weight9_20_2), .reg_activation12(reg_activation9_20_1), .reg_activation22(reg_activation9_20_2), .weight_en(weight_en));
SA22 U9_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_21_1), .partial_sum_in12(reg_psum8_21_2), .weight_in11(reg_weight8_21_1), .weight_in12(reg_weight8_21_2), .activation_in11(reg_activation9_20_1), .activation_in21(reg_activation9_20_2), .reg_partial_sum21(reg_psum9_21_1), .reg_partial_sum22(reg_psum9_21_2), .reg_weight21(reg_weight9_21_1), .reg_weight22(reg_weight9_21_2), .reg_activation12(reg_activation9_21_1), .reg_activation22(reg_activation9_21_2), .weight_en(weight_en));
SA22 U9_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_22_1), .partial_sum_in12(reg_psum8_22_2), .weight_in11(reg_weight8_22_1), .weight_in12(reg_weight8_22_2), .activation_in11(reg_activation9_21_1), .activation_in21(reg_activation9_21_2), .reg_partial_sum21(reg_psum9_22_1), .reg_partial_sum22(reg_psum9_22_2), .reg_weight21(reg_weight9_22_1), .reg_weight22(reg_weight9_22_2), .reg_activation12(reg_activation9_22_1), .reg_activation22(reg_activation9_22_2), .weight_en(weight_en));
SA22 U9_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_23_1), .partial_sum_in12(reg_psum8_23_2), .weight_in11(reg_weight8_23_1), .weight_in12(reg_weight8_23_2), .activation_in11(reg_activation9_22_1), .activation_in21(reg_activation9_22_2), .reg_partial_sum21(reg_psum9_23_1), .reg_partial_sum22(reg_psum9_23_2), .reg_weight21(reg_weight9_23_1), .reg_weight22(reg_weight9_23_2), .reg_activation12(reg_activation9_23_1), .reg_activation22(reg_activation9_23_2), .weight_en(weight_en));
SA22 U9_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_24_1), .partial_sum_in12(reg_psum8_24_2), .weight_in11(reg_weight8_24_1), .weight_in12(reg_weight8_24_2), .activation_in11(reg_activation9_23_1), .activation_in21(reg_activation9_23_2), .reg_partial_sum21(reg_psum9_24_1), .reg_partial_sum22(reg_psum9_24_2), .reg_weight21(reg_weight9_24_1), .reg_weight22(reg_weight9_24_2), .reg_activation12(reg_activation9_24_1), .reg_activation22(reg_activation9_24_2), .weight_en(weight_en));
SA22 U9_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_25_1), .partial_sum_in12(reg_psum8_25_2), .weight_in11(reg_weight8_25_1), .weight_in12(reg_weight8_25_2), .activation_in11(reg_activation9_24_1), .activation_in21(reg_activation9_24_2), .reg_partial_sum21(reg_psum9_25_1), .reg_partial_sum22(reg_psum9_25_2), .reg_weight21(reg_weight9_25_1), .reg_weight22(reg_weight9_25_2), .reg_activation12(reg_activation9_25_1), .reg_activation22(reg_activation9_25_2), .weight_en(weight_en));
SA22 U9_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_26_1), .partial_sum_in12(reg_psum8_26_2), .weight_in11(reg_weight8_26_1), .weight_in12(reg_weight8_26_2), .activation_in11(reg_activation9_25_1), .activation_in21(reg_activation9_25_2), .reg_partial_sum21(reg_psum9_26_1), .reg_partial_sum22(reg_psum9_26_2), .reg_weight21(reg_weight9_26_1), .reg_weight22(reg_weight9_26_2), .reg_activation12(reg_activation9_26_1), .reg_activation22(reg_activation9_26_2), .weight_en(weight_en));
SA22 U9_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_27_1), .partial_sum_in12(reg_psum8_27_2), .weight_in11(reg_weight8_27_1), .weight_in12(reg_weight8_27_2), .activation_in11(reg_activation9_26_1), .activation_in21(reg_activation9_26_2), .reg_partial_sum21(reg_psum9_27_1), .reg_partial_sum22(reg_psum9_27_2), .reg_weight21(reg_weight9_27_1), .reg_weight22(reg_weight9_27_2), .reg_activation12(reg_activation9_27_1), .reg_activation22(reg_activation9_27_2), .weight_en(weight_en));
SA22 U9_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_28_1), .partial_sum_in12(reg_psum8_28_2), .weight_in11(reg_weight8_28_1), .weight_in12(reg_weight8_28_2), .activation_in11(reg_activation9_27_1), .activation_in21(reg_activation9_27_2), .reg_partial_sum21(reg_psum9_28_1), .reg_partial_sum22(reg_psum9_28_2), .reg_weight21(reg_weight9_28_1), .reg_weight22(reg_weight9_28_2), .reg_activation12(reg_activation9_28_1), .reg_activation22(reg_activation9_28_2), .weight_en(weight_en));
SA22 U9_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_29_1), .partial_sum_in12(reg_psum8_29_2), .weight_in11(reg_weight8_29_1), .weight_in12(reg_weight8_29_2), .activation_in11(reg_activation9_28_1), .activation_in21(reg_activation9_28_2), .reg_partial_sum21(reg_psum9_29_1), .reg_partial_sum22(reg_psum9_29_2), .reg_weight21(reg_weight9_29_1), .reg_weight22(reg_weight9_29_2), .reg_activation12(reg_activation9_29_1), .reg_activation22(reg_activation9_29_2), .weight_en(weight_en));
SA22 U9_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_30_1), .partial_sum_in12(reg_psum8_30_2), .weight_in11(reg_weight8_30_1), .weight_in12(reg_weight8_30_2), .activation_in11(reg_activation9_29_1), .activation_in21(reg_activation9_29_2), .reg_partial_sum21(reg_psum9_30_1), .reg_partial_sum22(reg_psum9_30_2), .reg_weight21(reg_weight9_30_1), .reg_weight22(reg_weight9_30_2), .reg_activation12(reg_activation9_30_1), .reg_activation22(reg_activation9_30_2), .weight_en(weight_en));
SA22 U9_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_31_1), .partial_sum_in12(reg_psum8_31_2), .weight_in11(reg_weight8_31_1), .weight_in12(reg_weight8_31_2), .activation_in11(reg_activation9_30_1), .activation_in21(reg_activation9_30_2), .reg_partial_sum21(reg_psum9_31_1), .reg_partial_sum22(reg_psum9_31_2), .reg_weight21(reg_weight9_31_1), .reg_weight22(reg_weight9_31_2), .reg_activation12(reg_activation9_31_1), .reg_activation22(reg_activation9_31_2), .weight_en(weight_en));
SA22 U9_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum8_32_1), .partial_sum_in12(reg_psum8_32_2), .weight_in11(reg_weight8_32_1), .weight_in12(reg_weight8_32_2), .activation_in11(reg_activation9_31_1), .activation_in21(reg_activation9_31_2), .reg_partial_sum21(reg_psum9_32_1), .reg_partial_sum22(reg_psum9_32_2), .reg_weight21(reg_weight9_32_1), .reg_weight22(reg_weight9_32_2), .weight_en(weight_en));
SA22 U10_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_1_1), .partial_sum_in12(reg_psum9_1_2), .weight_in11(reg_weight9_1_1), .weight_in12(reg_weight9_1_2), .activation_in11(in_activation10_1_1), .activation_in21(in_activation10_1_2), .reg_partial_sum21(reg_psum10_1_1), .reg_partial_sum22(reg_psum10_1_2), .reg_weight21(reg_weight10_1_1), .reg_weight22(reg_weight10_1_2), .reg_activation12(reg_activation10_1_1), .reg_activation22(reg_activation10_1_2), .weight_en(weight_en));
SA22 U10_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_2_1), .partial_sum_in12(reg_psum9_2_2), .weight_in11(reg_weight9_2_1), .weight_in12(reg_weight9_2_2), .activation_in11(reg_activation10_1_1), .activation_in21(reg_activation10_1_2), .reg_partial_sum21(reg_psum10_2_1), .reg_partial_sum22(reg_psum10_2_2), .reg_weight21(reg_weight10_2_1), .reg_weight22(reg_weight10_2_2), .reg_activation12(reg_activation10_2_1), .reg_activation22(reg_activation10_2_2), .weight_en(weight_en));
SA22 U10_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_3_1), .partial_sum_in12(reg_psum9_3_2), .weight_in11(reg_weight9_3_1), .weight_in12(reg_weight9_3_2), .activation_in11(reg_activation10_2_1), .activation_in21(reg_activation10_2_2), .reg_partial_sum21(reg_psum10_3_1), .reg_partial_sum22(reg_psum10_3_2), .reg_weight21(reg_weight10_3_1), .reg_weight22(reg_weight10_3_2), .reg_activation12(reg_activation10_3_1), .reg_activation22(reg_activation10_3_2), .weight_en(weight_en));
SA22 U10_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_4_1), .partial_sum_in12(reg_psum9_4_2), .weight_in11(reg_weight9_4_1), .weight_in12(reg_weight9_4_2), .activation_in11(reg_activation10_3_1), .activation_in21(reg_activation10_3_2), .reg_partial_sum21(reg_psum10_4_1), .reg_partial_sum22(reg_psum10_4_2), .reg_weight21(reg_weight10_4_1), .reg_weight22(reg_weight10_4_2), .reg_activation12(reg_activation10_4_1), .reg_activation22(reg_activation10_4_2), .weight_en(weight_en));
SA22 U10_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_5_1), .partial_sum_in12(reg_psum9_5_2), .weight_in11(reg_weight9_5_1), .weight_in12(reg_weight9_5_2), .activation_in11(reg_activation10_4_1), .activation_in21(reg_activation10_4_2), .reg_partial_sum21(reg_psum10_5_1), .reg_partial_sum22(reg_psum10_5_2), .reg_weight21(reg_weight10_5_1), .reg_weight22(reg_weight10_5_2), .reg_activation12(reg_activation10_5_1), .reg_activation22(reg_activation10_5_2), .weight_en(weight_en));
SA22 U10_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_6_1), .partial_sum_in12(reg_psum9_6_2), .weight_in11(reg_weight9_6_1), .weight_in12(reg_weight9_6_2), .activation_in11(reg_activation10_5_1), .activation_in21(reg_activation10_5_2), .reg_partial_sum21(reg_psum10_6_1), .reg_partial_sum22(reg_psum10_6_2), .reg_weight21(reg_weight10_6_1), .reg_weight22(reg_weight10_6_2), .reg_activation12(reg_activation10_6_1), .reg_activation22(reg_activation10_6_2), .weight_en(weight_en));
SA22 U10_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_7_1), .partial_sum_in12(reg_psum9_7_2), .weight_in11(reg_weight9_7_1), .weight_in12(reg_weight9_7_2), .activation_in11(reg_activation10_6_1), .activation_in21(reg_activation10_6_2), .reg_partial_sum21(reg_psum10_7_1), .reg_partial_sum22(reg_psum10_7_2), .reg_weight21(reg_weight10_7_1), .reg_weight22(reg_weight10_7_2), .reg_activation12(reg_activation10_7_1), .reg_activation22(reg_activation10_7_2), .weight_en(weight_en));
SA22 U10_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_8_1), .partial_sum_in12(reg_psum9_8_2), .weight_in11(reg_weight9_8_1), .weight_in12(reg_weight9_8_2), .activation_in11(reg_activation10_7_1), .activation_in21(reg_activation10_7_2), .reg_partial_sum21(reg_psum10_8_1), .reg_partial_sum22(reg_psum10_8_2), .reg_weight21(reg_weight10_8_1), .reg_weight22(reg_weight10_8_2), .reg_activation12(reg_activation10_8_1), .reg_activation22(reg_activation10_8_2), .weight_en(weight_en));
SA22 U10_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_9_1), .partial_sum_in12(reg_psum9_9_2), .weight_in11(reg_weight9_9_1), .weight_in12(reg_weight9_9_2), .activation_in11(reg_activation10_8_1), .activation_in21(reg_activation10_8_2), .reg_partial_sum21(reg_psum10_9_1), .reg_partial_sum22(reg_psum10_9_2), .reg_weight21(reg_weight10_9_1), .reg_weight22(reg_weight10_9_2), .reg_activation12(reg_activation10_9_1), .reg_activation22(reg_activation10_9_2), .weight_en(weight_en));
SA22 U10_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_10_1), .partial_sum_in12(reg_psum9_10_2), .weight_in11(reg_weight9_10_1), .weight_in12(reg_weight9_10_2), .activation_in11(reg_activation10_9_1), .activation_in21(reg_activation10_9_2), .reg_partial_sum21(reg_psum10_10_1), .reg_partial_sum22(reg_psum10_10_2), .reg_weight21(reg_weight10_10_1), .reg_weight22(reg_weight10_10_2), .reg_activation12(reg_activation10_10_1), .reg_activation22(reg_activation10_10_2), .weight_en(weight_en));
SA22 U10_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_11_1), .partial_sum_in12(reg_psum9_11_2), .weight_in11(reg_weight9_11_1), .weight_in12(reg_weight9_11_2), .activation_in11(reg_activation10_10_1), .activation_in21(reg_activation10_10_2), .reg_partial_sum21(reg_psum10_11_1), .reg_partial_sum22(reg_psum10_11_2), .reg_weight21(reg_weight10_11_1), .reg_weight22(reg_weight10_11_2), .reg_activation12(reg_activation10_11_1), .reg_activation22(reg_activation10_11_2), .weight_en(weight_en));
SA22 U10_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_12_1), .partial_sum_in12(reg_psum9_12_2), .weight_in11(reg_weight9_12_1), .weight_in12(reg_weight9_12_2), .activation_in11(reg_activation10_11_1), .activation_in21(reg_activation10_11_2), .reg_partial_sum21(reg_psum10_12_1), .reg_partial_sum22(reg_psum10_12_2), .reg_weight21(reg_weight10_12_1), .reg_weight22(reg_weight10_12_2), .reg_activation12(reg_activation10_12_1), .reg_activation22(reg_activation10_12_2), .weight_en(weight_en));
SA22 U10_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_13_1), .partial_sum_in12(reg_psum9_13_2), .weight_in11(reg_weight9_13_1), .weight_in12(reg_weight9_13_2), .activation_in11(reg_activation10_12_1), .activation_in21(reg_activation10_12_2), .reg_partial_sum21(reg_psum10_13_1), .reg_partial_sum22(reg_psum10_13_2), .reg_weight21(reg_weight10_13_1), .reg_weight22(reg_weight10_13_2), .reg_activation12(reg_activation10_13_1), .reg_activation22(reg_activation10_13_2), .weight_en(weight_en));
SA22 U10_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_14_1), .partial_sum_in12(reg_psum9_14_2), .weight_in11(reg_weight9_14_1), .weight_in12(reg_weight9_14_2), .activation_in11(reg_activation10_13_1), .activation_in21(reg_activation10_13_2), .reg_partial_sum21(reg_psum10_14_1), .reg_partial_sum22(reg_psum10_14_2), .reg_weight21(reg_weight10_14_1), .reg_weight22(reg_weight10_14_2), .reg_activation12(reg_activation10_14_1), .reg_activation22(reg_activation10_14_2), .weight_en(weight_en));
SA22 U10_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_15_1), .partial_sum_in12(reg_psum9_15_2), .weight_in11(reg_weight9_15_1), .weight_in12(reg_weight9_15_2), .activation_in11(reg_activation10_14_1), .activation_in21(reg_activation10_14_2), .reg_partial_sum21(reg_psum10_15_1), .reg_partial_sum22(reg_psum10_15_2), .reg_weight21(reg_weight10_15_1), .reg_weight22(reg_weight10_15_2), .reg_activation12(reg_activation10_15_1), .reg_activation22(reg_activation10_15_2), .weight_en(weight_en));
SA22 U10_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_16_1), .partial_sum_in12(reg_psum9_16_2), .weight_in11(reg_weight9_16_1), .weight_in12(reg_weight9_16_2), .activation_in11(reg_activation10_15_1), .activation_in21(reg_activation10_15_2), .reg_partial_sum21(reg_psum10_16_1), .reg_partial_sum22(reg_psum10_16_2), .reg_weight21(reg_weight10_16_1), .reg_weight22(reg_weight10_16_2), .reg_activation12(reg_activation10_16_1), .reg_activation22(reg_activation10_16_2), .weight_en(weight_en));
SA22 U10_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_17_1), .partial_sum_in12(reg_psum9_17_2), .weight_in11(reg_weight9_17_1), .weight_in12(reg_weight9_17_2), .activation_in11(reg_activation10_16_1), .activation_in21(reg_activation10_16_2), .reg_partial_sum21(reg_psum10_17_1), .reg_partial_sum22(reg_psum10_17_2), .reg_weight21(reg_weight10_17_1), .reg_weight22(reg_weight10_17_2), .reg_activation12(reg_activation10_17_1), .reg_activation22(reg_activation10_17_2), .weight_en(weight_en));
SA22 U10_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_18_1), .partial_sum_in12(reg_psum9_18_2), .weight_in11(reg_weight9_18_1), .weight_in12(reg_weight9_18_2), .activation_in11(reg_activation10_17_1), .activation_in21(reg_activation10_17_2), .reg_partial_sum21(reg_psum10_18_1), .reg_partial_sum22(reg_psum10_18_2), .reg_weight21(reg_weight10_18_1), .reg_weight22(reg_weight10_18_2), .reg_activation12(reg_activation10_18_1), .reg_activation22(reg_activation10_18_2), .weight_en(weight_en));
SA22 U10_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_19_1), .partial_sum_in12(reg_psum9_19_2), .weight_in11(reg_weight9_19_1), .weight_in12(reg_weight9_19_2), .activation_in11(reg_activation10_18_1), .activation_in21(reg_activation10_18_2), .reg_partial_sum21(reg_psum10_19_1), .reg_partial_sum22(reg_psum10_19_2), .reg_weight21(reg_weight10_19_1), .reg_weight22(reg_weight10_19_2), .reg_activation12(reg_activation10_19_1), .reg_activation22(reg_activation10_19_2), .weight_en(weight_en));
SA22 U10_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_20_1), .partial_sum_in12(reg_psum9_20_2), .weight_in11(reg_weight9_20_1), .weight_in12(reg_weight9_20_2), .activation_in11(reg_activation10_19_1), .activation_in21(reg_activation10_19_2), .reg_partial_sum21(reg_psum10_20_1), .reg_partial_sum22(reg_psum10_20_2), .reg_weight21(reg_weight10_20_1), .reg_weight22(reg_weight10_20_2), .reg_activation12(reg_activation10_20_1), .reg_activation22(reg_activation10_20_2), .weight_en(weight_en));
SA22 U10_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_21_1), .partial_sum_in12(reg_psum9_21_2), .weight_in11(reg_weight9_21_1), .weight_in12(reg_weight9_21_2), .activation_in11(reg_activation10_20_1), .activation_in21(reg_activation10_20_2), .reg_partial_sum21(reg_psum10_21_1), .reg_partial_sum22(reg_psum10_21_2), .reg_weight21(reg_weight10_21_1), .reg_weight22(reg_weight10_21_2), .reg_activation12(reg_activation10_21_1), .reg_activation22(reg_activation10_21_2), .weight_en(weight_en));
SA22 U10_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_22_1), .partial_sum_in12(reg_psum9_22_2), .weight_in11(reg_weight9_22_1), .weight_in12(reg_weight9_22_2), .activation_in11(reg_activation10_21_1), .activation_in21(reg_activation10_21_2), .reg_partial_sum21(reg_psum10_22_1), .reg_partial_sum22(reg_psum10_22_2), .reg_weight21(reg_weight10_22_1), .reg_weight22(reg_weight10_22_2), .reg_activation12(reg_activation10_22_1), .reg_activation22(reg_activation10_22_2), .weight_en(weight_en));
SA22 U10_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_23_1), .partial_sum_in12(reg_psum9_23_2), .weight_in11(reg_weight9_23_1), .weight_in12(reg_weight9_23_2), .activation_in11(reg_activation10_22_1), .activation_in21(reg_activation10_22_2), .reg_partial_sum21(reg_psum10_23_1), .reg_partial_sum22(reg_psum10_23_2), .reg_weight21(reg_weight10_23_1), .reg_weight22(reg_weight10_23_2), .reg_activation12(reg_activation10_23_1), .reg_activation22(reg_activation10_23_2), .weight_en(weight_en));
SA22 U10_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_24_1), .partial_sum_in12(reg_psum9_24_2), .weight_in11(reg_weight9_24_1), .weight_in12(reg_weight9_24_2), .activation_in11(reg_activation10_23_1), .activation_in21(reg_activation10_23_2), .reg_partial_sum21(reg_psum10_24_1), .reg_partial_sum22(reg_psum10_24_2), .reg_weight21(reg_weight10_24_1), .reg_weight22(reg_weight10_24_2), .reg_activation12(reg_activation10_24_1), .reg_activation22(reg_activation10_24_2), .weight_en(weight_en));
SA22 U10_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_25_1), .partial_sum_in12(reg_psum9_25_2), .weight_in11(reg_weight9_25_1), .weight_in12(reg_weight9_25_2), .activation_in11(reg_activation10_24_1), .activation_in21(reg_activation10_24_2), .reg_partial_sum21(reg_psum10_25_1), .reg_partial_sum22(reg_psum10_25_2), .reg_weight21(reg_weight10_25_1), .reg_weight22(reg_weight10_25_2), .reg_activation12(reg_activation10_25_1), .reg_activation22(reg_activation10_25_2), .weight_en(weight_en));
SA22 U10_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_26_1), .partial_sum_in12(reg_psum9_26_2), .weight_in11(reg_weight9_26_1), .weight_in12(reg_weight9_26_2), .activation_in11(reg_activation10_25_1), .activation_in21(reg_activation10_25_2), .reg_partial_sum21(reg_psum10_26_1), .reg_partial_sum22(reg_psum10_26_2), .reg_weight21(reg_weight10_26_1), .reg_weight22(reg_weight10_26_2), .reg_activation12(reg_activation10_26_1), .reg_activation22(reg_activation10_26_2), .weight_en(weight_en));
SA22 U10_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_27_1), .partial_sum_in12(reg_psum9_27_2), .weight_in11(reg_weight9_27_1), .weight_in12(reg_weight9_27_2), .activation_in11(reg_activation10_26_1), .activation_in21(reg_activation10_26_2), .reg_partial_sum21(reg_psum10_27_1), .reg_partial_sum22(reg_psum10_27_2), .reg_weight21(reg_weight10_27_1), .reg_weight22(reg_weight10_27_2), .reg_activation12(reg_activation10_27_1), .reg_activation22(reg_activation10_27_2), .weight_en(weight_en));
SA22 U10_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_28_1), .partial_sum_in12(reg_psum9_28_2), .weight_in11(reg_weight9_28_1), .weight_in12(reg_weight9_28_2), .activation_in11(reg_activation10_27_1), .activation_in21(reg_activation10_27_2), .reg_partial_sum21(reg_psum10_28_1), .reg_partial_sum22(reg_psum10_28_2), .reg_weight21(reg_weight10_28_1), .reg_weight22(reg_weight10_28_2), .reg_activation12(reg_activation10_28_1), .reg_activation22(reg_activation10_28_2), .weight_en(weight_en));
SA22 U10_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_29_1), .partial_sum_in12(reg_psum9_29_2), .weight_in11(reg_weight9_29_1), .weight_in12(reg_weight9_29_2), .activation_in11(reg_activation10_28_1), .activation_in21(reg_activation10_28_2), .reg_partial_sum21(reg_psum10_29_1), .reg_partial_sum22(reg_psum10_29_2), .reg_weight21(reg_weight10_29_1), .reg_weight22(reg_weight10_29_2), .reg_activation12(reg_activation10_29_1), .reg_activation22(reg_activation10_29_2), .weight_en(weight_en));
SA22 U10_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_30_1), .partial_sum_in12(reg_psum9_30_2), .weight_in11(reg_weight9_30_1), .weight_in12(reg_weight9_30_2), .activation_in11(reg_activation10_29_1), .activation_in21(reg_activation10_29_2), .reg_partial_sum21(reg_psum10_30_1), .reg_partial_sum22(reg_psum10_30_2), .reg_weight21(reg_weight10_30_1), .reg_weight22(reg_weight10_30_2), .reg_activation12(reg_activation10_30_1), .reg_activation22(reg_activation10_30_2), .weight_en(weight_en));
SA22 U10_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_31_1), .partial_sum_in12(reg_psum9_31_2), .weight_in11(reg_weight9_31_1), .weight_in12(reg_weight9_31_2), .activation_in11(reg_activation10_30_1), .activation_in21(reg_activation10_30_2), .reg_partial_sum21(reg_psum10_31_1), .reg_partial_sum22(reg_psum10_31_2), .reg_weight21(reg_weight10_31_1), .reg_weight22(reg_weight10_31_2), .reg_activation12(reg_activation10_31_1), .reg_activation22(reg_activation10_31_2), .weight_en(weight_en));
SA22 U10_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum9_32_1), .partial_sum_in12(reg_psum9_32_2), .weight_in11(reg_weight9_32_1), .weight_in12(reg_weight9_32_2), .activation_in11(reg_activation10_31_1), .activation_in21(reg_activation10_31_2), .reg_partial_sum21(reg_psum10_32_1), .reg_partial_sum22(reg_psum10_32_2), .reg_weight21(reg_weight10_32_1), .reg_weight22(reg_weight10_32_2), .weight_en(weight_en));
SA22 U11_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_1_1), .partial_sum_in12(reg_psum10_1_2), .weight_in11(reg_weight10_1_1), .weight_in12(reg_weight10_1_2), .activation_in11(in_activation11_1_1), .activation_in21(in_activation11_1_2), .reg_partial_sum21(reg_psum11_1_1), .reg_partial_sum22(reg_psum11_1_2), .reg_weight21(reg_weight11_1_1), .reg_weight22(reg_weight11_1_2), .reg_activation12(reg_activation11_1_1), .reg_activation22(reg_activation11_1_2), .weight_en(weight_en));
SA22 U11_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_2_1), .partial_sum_in12(reg_psum10_2_2), .weight_in11(reg_weight10_2_1), .weight_in12(reg_weight10_2_2), .activation_in11(reg_activation11_1_1), .activation_in21(reg_activation11_1_2), .reg_partial_sum21(reg_psum11_2_1), .reg_partial_sum22(reg_psum11_2_2), .reg_weight21(reg_weight11_2_1), .reg_weight22(reg_weight11_2_2), .reg_activation12(reg_activation11_2_1), .reg_activation22(reg_activation11_2_2), .weight_en(weight_en));
SA22 U11_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_3_1), .partial_sum_in12(reg_psum10_3_2), .weight_in11(reg_weight10_3_1), .weight_in12(reg_weight10_3_2), .activation_in11(reg_activation11_2_1), .activation_in21(reg_activation11_2_2), .reg_partial_sum21(reg_psum11_3_1), .reg_partial_sum22(reg_psum11_3_2), .reg_weight21(reg_weight11_3_1), .reg_weight22(reg_weight11_3_2), .reg_activation12(reg_activation11_3_1), .reg_activation22(reg_activation11_3_2), .weight_en(weight_en));
SA22 U11_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_4_1), .partial_sum_in12(reg_psum10_4_2), .weight_in11(reg_weight10_4_1), .weight_in12(reg_weight10_4_2), .activation_in11(reg_activation11_3_1), .activation_in21(reg_activation11_3_2), .reg_partial_sum21(reg_psum11_4_1), .reg_partial_sum22(reg_psum11_4_2), .reg_weight21(reg_weight11_4_1), .reg_weight22(reg_weight11_4_2), .reg_activation12(reg_activation11_4_1), .reg_activation22(reg_activation11_4_2), .weight_en(weight_en));
SA22 U11_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_5_1), .partial_sum_in12(reg_psum10_5_2), .weight_in11(reg_weight10_5_1), .weight_in12(reg_weight10_5_2), .activation_in11(reg_activation11_4_1), .activation_in21(reg_activation11_4_2), .reg_partial_sum21(reg_psum11_5_1), .reg_partial_sum22(reg_psum11_5_2), .reg_weight21(reg_weight11_5_1), .reg_weight22(reg_weight11_5_2), .reg_activation12(reg_activation11_5_1), .reg_activation22(reg_activation11_5_2), .weight_en(weight_en));
SA22 U11_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_6_1), .partial_sum_in12(reg_psum10_6_2), .weight_in11(reg_weight10_6_1), .weight_in12(reg_weight10_6_2), .activation_in11(reg_activation11_5_1), .activation_in21(reg_activation11_5_2), .reg_partial_sum21(reg_psum11_6_1), .reg_partial_sum22(reg_psum11_6_2), .reg_weight21(reg_weight11_6_1), .reg_weight22(reg_weight11_6_2), .reg_activation12(reg_activation11_6_1), .reg_activation22(reg_activation11_6_2), .weight_en(weight_en));
SA22 U11_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_7_1), .partial_sum_in12(reg_psum10_7_2), .weight_in11(reg_weight10_7_1), .weight_in12(reg_weight10_7_2), .activation_in11(reg_activation11_6_1), .activation_in21(reg_activation11_6_2), .reg_partial_sum21(reg_psum11_7_1), .reg_partial_sum22(reg_psum11_7_2), .reg_weight21(reg_weight11_7_1), .reg_weight22(reg_weight11_7_2), .reg_activation12(reg_activation11_7_1), .reg_activation22(reg_activation11_7_2), .weight_en(weight_en));
SA22 U11_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_8_1), .partial_sum_in12(reg_psum10_8_2), .weight_in11(reg_weight10_8_1), .weight_in12(reg_weight10_8_2), .activation_in11(reg_activation11_7_1), .activation_in21(reg_activation11_7_2), .reg_partial_sum21(reg_psum11_8_1), .reg_partial_sum22(reg_psum11_8_2), .reg_weight21(reg_weight11_8_1), .reg_weight22(reg_weight11_8_2), .reg_activation12(reg_activation11_8_1), .reg_activation22(reg_activation11_8_2), .weight_en(weight_en));
SA22 U11_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_9_1), .partial_sum_in12(reg_psum10_9_2), .weight_in11(reg_weight10_9_1), .weight_in12(reg_weight10_9_2), .activation_in11(reg_activation11_8_1), .activation_in21(reg_activation11_8_2), .reg_partial_sum21(reg_psum11_9_1), .reg_partial_sum22(reg_psum11_9_2), .reg_weight21(reg_weight11_9_1), .reg_weight22(reg_weight11_9_2), .reg_activation12(reg_activation11_9_1), .reg_activation22(reg_activation11_9_2), .weight_en(weight_en));
SA22 U11_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_10_1), .partial_sum_in12(reg_psum10_10_2), .weight_in11(reg_weight10_10_1), .weight_in12(reg_weight10_10_2), .activation_in11(reg_activation11_9_1), .activation_in21(reg_activation11_9_2), .reg_partial_sum21(reg_psum11_10_1), .reg_partial_sum22(reg_psum11_10_2), .reg_weight21(reg_weight11_10_1), .reg_weight22(reg_weight11_10_2), .reg_activation12(reg_activation11_10_1), .reg_activation22(reg_activation11_10_2), .weight_en(weight_en));
SA22 U11_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_11_1), .partial_sum_in12(reg_psum10_11_2), .weight_in11(reg_weight10_11_1), .weight_in12(reg_weight10_11_2), .activation_in11(reg_activation11_10_1), .activation_in21(reg_activation11_10_2), .reg_partial_sum21(reg_psum11_11_1), .reg_partial_sum22(reg_psum11_11_2), .reg_weight21(reg_weight11_11_1), .reg_weight22(reg_weight11_11_2), .reg_activation12(reg_activation11_11_1), .reg_activation22(reg_activation11_11_2), .weight_en(weight_en));
SA22 U11_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_12_1), .partial_sum_in12(reg_psum10_12_2), .weight_in11(reg_weight10_12_1), .weight_in12(reg_weight10_12_2), .activation_in11(reg_activation11_11_1), .activation_in21(reg_activation11_11_2), .reg_partial_sum21(reg_psum11_12_1), .reg_partial_sum22(reg_psum11_12_2), .reg_weight21(reg_weight11_12_1), .reg_weight22(reg_weight11_12_2), .reg_activation12(reg_activation11_12_1), .reg_activation22(reg_activation11_12_2), .weight_en(weight_en));
SA22 U11_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_13_1), .partial_sum_in12(reg_psum10_13_2), .weight_in11(reg_weight10_13_1), .weight_in12(reg_weight10_13_2), .activation_in11(reg_activation11_12_1), .activation_in21(reg_activation11_12_2), .reg_partial_sum21(reg_psum11_13_1), .reg_partial_sum22(reg_psum11_13_2), .reg_weight21(reg_weight11_13_1), .reg_weight22(reg_weight11_13_2), .reg_activation12(reg_activation11_13_1), .reg_activation22(reg_activation11_13_2), .weight_en(weight_en));
SA22 U11_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_14_1), .partial_sum_in12(reg_psum10_14_2), .weight_in11(reg_weight10_14_1), .weight_in12(reg_weight10_14_2), .activation_in11(reg_activation11_13_1), .activation_in21(reg_activation11_13_2), .reg_partial_sum21(reg_psum11_14_1), .reg_partial_sum22(reg_psum11_14_2), .reg_weight21(reg_weight11_14_1), .reg_weight22(reg_weight11_14_2), .reg_activation12(reg_activation11_14_1), .reg_activation22(reg_activation11_14_2), .weight_en(weight_en));
SA22 U11_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_15_1), .partial_sum_in12(reg_psum10_15_2), .weight_in11(reg_weight10_15_1), .weight_in12(reg_weight10_15_2), .activation_in11(reg_activation11_14_1), .activation_in21(reg_activation11_14_2), .reg_partial_sum21(reg_psum11_15_1), .reg_partial_sum22(reg_psum11_15_2), .reg_weight21(reg_weight11_15_1), .reg_weight22(reg_weight11_15_2), .reg_activation12(reg_activation11_15_1), .reg_activation22(reg_activation11_15_2), .weight_en(weight_en));
SA22 U11_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_16_1), .partial_sum_in12(reg_psum10_16_2), .weight_in11(reg_weight10_16_1), .weight_in12(reg_weight10_16_2), .activation_in11(reg_activation11_15_1), .activation_in21(reg_activation11_15_2), .reg_partial_sum21(reg_psum11_16_1), .reg_partial_sum22(reg_psum11_16_2), .reg_weight21(reg_weight11_16_1), .reg_weight22(reg_weight11_16_2), .reg_activation12(reg_activation11_16_1), .reg_activation22(reg_activation11_16_2), .weight_en(weight_en));
SA22 U11_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_17_1), .partial_sum_in12(reg_psum10_17_2), .weight_in11(reg_weight10_17_1), .weight_in12(reg_weight10_17_2), .activation_in11(reg_activation11_16_1), .activation_in21(reg_activation11_16_2), .reg_partial_sum21(reg_psum11_17_1), .reg_partial_sum22(reg_psum11_17_2), .reg_weight21(reg_weight11_17_1), .reg_weight22(reg_weight11_17_2), .reg_activation12(reg_activation11_17_1), .reg_activation22(reg_activation11_17_2), .weight_en(weight_en));
SA22 U11_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_18_1), .partial_sum_in12(reg_psum10_18_2), .weight_in11(reg_weight10_18_1), .weight_in12(reg_weight10_18_2), .activation_in11(reg_activation11_17_1), .activation_in21(reg_activation11_17_2), .reg_partial_sum21(reg_psum11_18_1), .reg_partial_sum22(reg_psum11_18_2), .reg_weight21(reg_weight11_18_1), .reg_weight22(reg_weight11_18_2), .reg_activation12(reg_activation11_18_1), .reg_activation22(reg_activation11_18_2), .weight_en(weight_en));
SA22 U11_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_19_1), .partial_sum_in12(reg_psum10_19_2), .weight_in11(reg_weight10_19_1), .weight_in12(reg_weight10_19_2), .activation_in11(reg_activation11_18_1), .activation_in21(reg_activation11_18_2), .reg_partial_sum21(reg_psum11_19_1), .reg_partial_sum22(reg_psum11_19_2), .reg_weight21(reg_weight11_19_1), .reg_weight22(reg_weight11_19_2), .reg_activation12(reg_activation11_19_1), .reg_activation22(reg_activation11_19_2), .weight_en(weight_en));
SA22 U11_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_20_1), .partial_sum_in12(reg_psum10_20_2), .weight_in11(reg_weight10_20_1), .weight_in12(reg_weight10_20_2), .activation_in11(reg_activation11_19_1), .activation_in21(reg_activation11_19_2), .reg_partial_sum21(reg_psum11_20_1), .reg_partial_sum22(reg_psum11_20_2), .reg_weight21(reg_weight11_20_1), .reg_weight22(reg_weight11_20_2), .reg_activation12(reg_activation11_20_1), .reg_activation22(reg_activation11_20_2), .weight_en(weight_en));
SA22 U11_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_21_1), .partial_sum_in12(reg_psum10_21_2), .weight_in11(reg_weight10_21_1), .weight_in12(reg_weight10_21_2), .activation_in11(reg_activation11_20_1), .activation_in21(reg_activation11_20_2), .reg_partial_sum21(reg_psum11_21_1), .reg_partial_sum22(reg_psum11_21_2), .reg_weight21(reg_weight11_21_1), .reg_weight22(reg_weight11_21_2), .reg_activation12(reg_activation11_21_1), .reg_activation22(reg_activation11_21_2), .weight_en(weight_en));
SA22 U11_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_22_1), .partial_sum_in12(reg_psum10_22_2), .weight_in11(reg_weight10_22_1), .weight_in12(reg_weight10_22_2), .activation_in11(reg_activation11_21_1), .activation_in21(reg_activation11_21_2), .reg_partial_sum21(reg_psum11_22_1), .reg_partial_sum22(reg_psum11_22_2), .reg_weight21(reg_weight11_22_1), .reg_weight22(reg_weight11_22_2), .reg_activation12(reg_activation11_22_1), .reg_activation22(reg_activation11_22_2), .weight_en(weight_en));
SA22 U11_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_23_1), .partial_sum_in12(reg_psum10_23_2), .weight_in11(reg_weight10_23_1), .weight_in12(reg_weight10_23_2), .activation_in11(reg_activation11_22_1), .activation_in21(reg_activation11_22_2), .reg_partial_sum21(reg_psum11_23_1), .reg_partial_sum22(reg_psum11_23_2), .reg_weight21(reg_weight11_23_1), .reg_weight22(reg_weight11_23_2), .reg_activation12(reg_activation11_23_1), .reg_activation22(reg_activation11_23_2), .weight_en(weight_en));
SA22 U11_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_24_1), .partial_sum_in12(reg_psum10_24_2), .weight_in11(reg_weight10_24_1), .weight_in12(reg_weight10_24_2), .activation_in11(reg_activation11_23_1), .activation_in21(reg_activation11_23_2), .reg_partial_sum21(reg_psum11_24_1), .reg_partial_sum22(reg_psum11_24_2), .reg_weight21(reg_weight11_24_1), .reg_weight22(reg_weight11_24_2), .reg_activation12(reg_activation11_24_1), .reg_activation22(reg_activation11_24_2), .weight_en(weight_en));
SA22 U11_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_25_1), .partial_sum_in12(reg_psum10_25_2), .weight_in11(reg_weight10_25_1), .weight_in12(reg_weight10_25_2), .activation_in11(reg_activation11_24_1), .activation_in21(reg_activation11_24_2), .reg_partial_sum21(reg_psum11_25_1), .reg_partial_sum22(reg_psum11_25_2), .reg_weight21(reg_weight11_25_1), .reg_weight22(reg_weight11_25_2), .reg_activation12(reg_activation11_25_1), .reg_activation22(reg_activation11_25_2), .weight_en(weight_en));
SA22 U11_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_26_1), .partial_sum_in12(reg_psum10_26_2), .weight_in11(reg_weight10_26_1), .weight_in12(reg_weight10_26_2), .activation_in11(reg_activation11_25_1), .activation_in21(reg_activation11_25_2), .reg_partial_sum21(reg_psum11_26_1), .reg_partial_sum22(reg_psum11_26_2), .reg_weight21(reg_weight11_26_1), .reg_weight22(reg_weight11_26_2), .reg_activation12(reg_activation11_26_1), .reg_activation22(reg_activation11_26_2), .weight_en(weight_en));
SA22 U11_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_27_1), .partial_sum_in12(reg_psum10_27_2), .weight_in11(reg_weight10_27_1), .weight_in12(reg_weight10_27_2), .activation_in11(reg_activation11_26_1), .activation_in21(reg_activation11_26_2), .reg_partial_sum21(reg_psum11_27_1), .reg_partial_sum22(reg_psum11_27_2), .reg_weight21(reg_weight11_27_1), .reg_weight22(reg_weight11_27_2), .reg_activation12(reg_activation11_27_1), .reg_activation22(reg_activation11_27_2), .weight_en(weight_en));
SA22 U11_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_28_1), .partial_sum_in12(reg_psum10_28_2), .weight_in11(reg_weight10_28_1), .weight_in12(reg_weight10_28_2), .activation_in11(reg_activation11_27_1), .activation_in21(reg_activation11_27_2), .reg_partial_sum21(reg_psum11_28_1), .reg_partial_sum22(reg_psum11_28_2), .reg_weight21(reg_weight11_28_1), .reg_weight22(reg_weight11_28_2), .reg_activation12(reg_activation11_28_1), .reg_activation22(reg_activation11_28_2), .weight_en(weight_en));
SA22 U11_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_29_1), .partial_sum_in12(reg_psum10_29_2), .weight_in11(reg_weight10_29_1), .weight_in12(reg_weight10_29_2), .activation_in11(reg_activation11_28_1), .activation_in21(reg_activation11_28_2), .reg_partial_sum21(reg_psum11_29_1), .reg_partial_sum22(reg_psum11_29_2), .reg_weight21(reg_weight11_29_1), .reg_weight22(reg_weight11_29_2), .reg_activation12(reg_activation11_29_1), .reg_activation22(reg_activation11_29_2), .weight_en(weight_en));
SA22 U11_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_30_1), .partial_sum_in12(reg_psum10_30_2), .weight_in11(reg_weight10_30_1), .weight_in12(reg_weight10_30_2), .activation_in11(reg_activation11_29_1), .activation_in21(reg_activation11_29_2), .reg_partial_sum21(reg_psum11_30_1), .reg_partial_sum22(reg_psum11_30_2), .reg_weight21(reg_weight11_30_1), .reg_weight22(reg_weight11_30_2), .reg_activation12(reg_activation11_30_1), .reg_activation22(reg_activation11_30_2), .weight_en(weight_en));
SA22 U11_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_31_1), .partial_sum_in12(reg_psum10_31_2), .weight_in11(reg_weight10_31_1), .weight_in12(reg_weight10_31_2), .activation_in11(reg_activation11_30_1), .activation_in21(reg_activation11_30_2), .reg_partial_sum21(reg_psum11_31_1), .reg_partial_sum22(reg_psum11_31_2), .reg_weight21(reg_weight11_31_1), .reg_weight22(reg_weight11_31_2), .reg_activation12(reg_activation11_31_1), .reg_activation22(reg_activation11_31_2), .weight_en(weight_en));
SA22 U11_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum10_32_1), .partial_sum_in12(reg_psum10_32_2), .weight_in11(reg_weight10_32_1), .weight_in12(reg_weight10_32_2), .activation_in11(reg_activation11_31_1), .activation_in21(reg_activation11_31_2), .reg_partial_sum21(reg_psum11_32_1), .reg_partial_sum22(reg_psum11_32_2), .reg_weight21(reg_weight11_32_1), .reg_weight22(reg_weight11_32_2), .weight_en(weight_en));
SA22 U12_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_1_1), .partial_sum_in12(reg_psum11_1_2), .weight_in11(reg_weight11_1_1), .weight_in12(reg_weight11_1_2), .activation_in11(in_activation12_1_1), .activation_in21(in_activation12_1_2), .reg_partial_sum21(reg_psum12_1_1), .reg_partial_sum22(reg_psum12_1_2), .reg_weight21(reg_weight12_1_1), .reg_weight22(reg_weight12_1_2), .reg_activation12(reg_activation12_1_1), .reg_activation22(reg_activation12_1_2), .weight_en(weight_en));
SA22 U12_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_2_1), .partial_sum_in12(reg_psum11_2_2), .weight_in11(reg_weight11_2_1), .weight_in12(reg_weight11_2_2), .activation_in11(reg_activation12_1_1), .activation_in21(reg_activation12_1_2), .reg_partial_sum21(reg_psum12_2_1), .reg_partial_sum22(reg_psum12_2_2), .reg_weight21(reg_weight12_2_1), .reg_weight22(reg_weight12_2_2), .reg_activation12(reg_activation12_2_1), .reg_activation22(reg_activation12_2_2), .weight_en(weight_en));
SA22 U12_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_3_1), .partial_sum_in12(reg_psum11_3_2), .weight_in11(reg_weight11_3_1), .weight_in12(reg_weight11_3_2), .activation_in11(reg_activation12_2_1), .activation_in21(reg_activation12_2_2), .reg_partial_sum21(reg_psum12_3_1), .reg_partial_sum22(reg_psum12_3_2), .reg_weight21(reg_weight12_3_1), .reg_weight22(reg_weight12_3_2), .reg_activation12(reg_activation12_3_1), .reg_activation22(reg_activation12_3_2), .weight_en(weight_en));
SA22 U12_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_4_1), .partial_sum_in12(reg_psum11_4_2), .weight_in11(reg_weight11_4_1), .weight_in12(reg_weight11_4_2), .activation_in11(reg_activation12_3_1), .activation_in21(reg_activation12_3_2), .reg_partial_sum21(reg_psum12_4_1), .reg_partial_sum22(reg_psum12_4_2), .reg_weight21(reg_weight12_4_1), .reg_weight22(reg_weight12_4_2), .reg_activation12(reg_activation12_4_1), .reg_activation22(reg_activation12_4_2), .weight_en(weight_en));
SA22 U12_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_5_1), .partial_sum_in12(reg_psum11_5_2), .weight_in11(reg_weight11_5_1), .weight_in12(reg_weight11_5_2), .activation_in11(reg_activation12_4_1), .activation_in21(reg_activation12_4_2), .reg_partial_sum21(reg_psum12_5_1), .reg_partial_sum22(reg_psum12_5_2), .reg_weight21(reg_weight12_5_1), .reg_weight22(reg_weight12_5_2), .reg_activation12(reg_activation12_5_1), .reg_activation22(reg_activation12_5_2), .weight_en(weight_en));
SA22 U12_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_6_1), .partial_sum_in12(reg_psum11_6_2), .weight_in11(reg_weight11_6_1), .weight_in12(reg_weight11_6_2), .activation_in11(reg_activation12_5_1), .activation_in21(reg_activation12_5_2), .reg_partial_sum21(reg_psum12_6_1), .reg_partial_sum22(reg_psum12_6_2), .reg_weight21(reg_weight12_6_1), .reg_weight22(reg_weight12_6_2), .reg_activation12(reg_activation12_6_1), .reg_activation22(reg_activation12_6_2), .weight_en(weight_en));
SA22 U12_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_7_1), .partial_sum_in12(reg_psum11_7_2), .weight_in11(reg_weight11_7_1), .weight_in12(reg_weight11_7_2), .activation_in11(reg_activation12_6_1), .activation_in21(reg_activation12_6_2), .reg_partial_sum21(reg_psum12_7_1), .reg_partial_sum22(reg_psum12_7_2), .reg_weight21(reg_weight12_7_1), .reg_weight22(reg_weight12_7_2), .reg_activation12(reg_activation12_7_1), .reg_activation22(reg_activation12_7_2), .weight_en(weight_en));
SA22 U12_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_8_1), .partial_sum_in12(reg_psum11_8_2), .weight_in11(reg_weight11_8_1), .weight_in12(reg_weight11_8_2), .activation_in11(reg_activation12_7_1), .activation_in21(reg_activation12_7_2), .reg_partial_sum21(reg_psum12_8_1), .reg_partial_sum22(reg_psum12_8_2), .reg_weight21(reg_weight12_8_1), .reg_weight22(reg_weight12_8_2), .reg_activation12(reg_activation12_8_1), .reg_activation22(reg_activation12_8_2), .weight_en(weight_en));
SA22 U12_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_9_1), .partial_sum_in12(reg_psum11_9_2), .weight_in11(reg_weight11_9_1), .weight_in12(reg_weight11_9_2), .activation_in11(reg_activation12_8_1), .activation_in21(reg_activation12_8_2), .reg_partial_sum21(reg_psum12_9_1), .reg_partial_sum22(reg_psum12_9_2), .reg_weight21(reg_weight12_9_1), .reg_weight22(reg_weight12_9_2), .reg_activation12(reg_activation12_9_1), .reg_activation22(reg_activation12_9_2), .weight_en(weight_en));
SA22 U12_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_10_1), .partial_sum_in12(reg_psum11_10_2), .weight_in11(reg_weight11_10_1), .weight_in12(reg_weight11_10_2), .activation_in11(reg_activation12_9_1), .activation_in21(reg_activation12_9_2), .reg_partial_sum21(reg_psum12_10_1), .reg_partial_sum22(reg_psum12_10_2), .reg_weight21(reg_weight12_10_1), .reg_weight22(reg_weight12_10_2), .reg_activation12(reg_activation12_10_1), .reg_activation22(reg_activation12_10_2), .weight_en(weight_en));
SA22 U12_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_11_1), .partial_sum_in12(reg_psum11_11_2), .weight_in11(reg_weight11_11_1), .weight_in12(reg_weight11_11_2), .activation_in11(reg_activation12_10_1), .activation_in21(reg_activation12_10_2), .reg_partial_sum21(reg_psum12_11_1), .reg_partial_sum22(reg_psum12_11_2), .reg_weight21(reg_weight12_11_1), .reg_weight22(reg_weight12_11_2), .reg_activation12(reg_activation12_11_1), .reg_activation22(reg_activation12_11_2), .weight_en(weight_en));
SA22 U12_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_12_1), .partial_sum_in12(reg_psum11_12_2), .weight_in11(reg_weight11_12_1), .weight_in12(reg_weight11_12_2), .activation_in11(reg_activation12_11_1), .activation_in21(reg_activation12_11_2), .reg_partial_sum21(reg_psum12_12_1), .reg_partial_sum22(reg_psum12_12_2), .reg_weight21(reg_weight12_12_1), .reg_weight22(reg_weight12_12_2), .reg_activation12(reg_activation12_12_1), .reg_activation22(reg_activation12_12_2), .weight_en(weight_en));
SA22 U12_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_13_1), .partial_sum_in12(reg_psum11_13_2), .weight_in11(reg_weight11_13_1), .weight_in12(reg_weight11_13_2), .activation_in11(reg_activation12_12_1), .activation_in21(reg_activation12_12_2), .reg_partial_sum21(reg_psum12_13_1), .reg_partial_sum22(reg_psum12_13_2), .reg_weight21(reg_weight12_13_1), .reg_weight22(reg_weight12_13_2), .reg_activation12(reg_activation12_13_1), .reg_activation22(reg_activation12_13_2), .weight_en(weight_en));
SA22 U12_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_14_1), .partial_sum_in12(reg_psum11_14_2), .weight_in11(reg_weight11_14_1), .weight_in12(reg_weight11_14_2), .activation_in11(reg_activation12_13_1), .activation_in21(reg_activation12_13_2), .reg_partial_sum21(reg_psum12_14_1), .reg_partial_sum22(reg_psum12_14_2), .reg_weight21(reg_weight12_14_1), .reg_weight22(reg_weight12_14_2), .reg_activation12(reg_activation12_14_1), .reg_activation22(reg_activation12_14_2), .weight_en(weight_en));
SA22 U12_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_15_1), .partial_sum_in12(reg_psum11_15_2), .weight_in11(reg_weight11_15_1), .weight_in12(reg_weight11_15_2), .activation_in11(reg_activation12_14_1), .activation_in21(reg_activation12_14_2), .reg_partial_sum21(reg_psum12_15_1), .reg_partial_sum22(reg_psum12_15_2), .reg_weight21(reg_weight12_15_1), .reg_weight22(reg_weight12_15_2), .reg_activation12(reg_activation12_15_1), .reg_activation22(reg_activation12_15_2), .weight_en(weight_en));
SA22 U12_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_16_1), .partial_sum_in12(reg_psum11_16_2), .weight_in11(reg_weight11_16_1), .weight_in12(reg_weight11_16_2), .activation_in11(reg_activation12_15_1), .activation_in21(reg_activation12_15_2), .reg_partial_sum21(reg_psum12_16_1), .reg_partial_sum22(reg_psum12_16_2), .reg_weight21(reg_weight12_16_1), .reg_weight22(reg_weight12_16_2), .reg_activation12(reg_activation12_16_1), .reg_activation22(reg_activation12_16_2), .weight_en(weight_en));
SA22 U12_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_17_1), .partial_sum_in12(reg_psum11_17_2), .weight_in11(reg_weight11_17_1), .weight_in12(reg_weight11_17_2), .activation_in11(reg_activation12_16_1), .activation_in21(reg_activation12_16_2), .reg_partial_sum21(reg_psum12_17_1), .reg_partial_sum22(reg_psum12_17_2), .reg_weight21(reg_weight12_17_1), .reg_weight22(reg_weight12_17_2), .reg_activation12(reg_activation12_17_1), .reg_activation22(reg_activation12_17_2), .weight_en(weight_en));
SA22 U12_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_18_1), .partial_sum_in12(reg_psum11_18_2), .weight_in11(reg_weight11_18_1), .weight_in12(reg_weight11_18_2), .activation_in11(reg_activation12_17_1), .activation_in21(reg_activation12_17_2), .reg_partial_sum21(reg_psum12_18_1), .reg_partial_sum22(reg_psum12_18_2), .reg_weight21(reg_weight12_18_1), .reg_weight22(reg_weight12_18_2), .reg_activation12(reg_activation12_18_1), .reg_activation22(reg_activation12_18_2), .weight_en(weight_en));
SA22 U12_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_19_1), .partial_sum_in12(reg_psum11_19_2), .weight_in11(reg_weight11_19_1), .weight_in12(reg_weight11_19_2), .activation_in11(reg_activation12_18_1), .activation_in21(reg_activation12_18_2), .reg_partial_sum21(reg_psum12_19_1), .reg_partial_sum22(reg_psum12_19_2), .reg_weight21(reg_weight12_19_1), .reg_weight22(reg_weight12_19_2), .reg_activation12(reg_activation12_19_1), .reg_activation22(reg_activation12_19_2), .weight_en(weight_en));
SA22 U12_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_20_1), .partial_sum_in12(reg_psum11_20_2), .weight_in11(reg_weight11_20_1), .weight_in12(reg_weight11_20_2), .activation_in11(reg_activation12_19_1), .activation_in21(reg_activation12_19_2), .reg_partial_sum21(reg_psum12_20_1), .reg_partial_sum22(reg_psum12_20_2), .reg_weight21(reg_weight12_20_1), .reg_weight22(reg_weight12_20_2), .reg_activation12(reg_activation12_20_1), .reg_activation22(reg_activation12_20_2), .weight_en(weight_en));
SA22 U12_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_21_1), .partial_sum_in12(reg_psum11_21_2), .weight_in11(reg_weight11_21_1), .weight_in12(reg_weight11_21_2), .activation_in11(reg_activation12_20_1), .activation_in21(reg_activation12_20_2), .reg_partial_sum21(reg_psum12_21_1), .reg_partial_sum22(reg_psum12_21_2), .reg_weight21(reg_weight12_21_1), .reg_weight22(reg_weight12_21_2), .reg_activation12(reg_activation12_21_1), .reg_activation22(reg_activation12_21_2), .weight_en(weight_en));
SA22 U12_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_22_1), .partial_sum_in12(reg_psum11_22_2), .weight_in11(reg_weight11_22_1), .weight_in12(reg_weight11_22_2), .activation_in11(reg_activation12_21_1), .activation_in21(reg_activation12_21_2), .reg_partial_sum21(reg_psum12_22_1), .reg_partial_sum22(reg_psum12_22_2), .reg_weight21(reg_weight12_22_1), .reg_weight22(reg_weight12_22_2), .reg_activation12(reg_activation12_22_1), .reg_activation22(reg_activation12_22_2), .weight_en(weight_en));
SA22 U12_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_23_1), .partial_sum_in12(reg_psum11_23_2), .weight_in11(reg_weight11_23_1), .weight_in12(reg_weight11_23_2), .activation_in11(reg_activation12_22_1), .activation_in21(reg_activation12_22_2), .reg_partial_sum21(reg_psum12_23_1), .reg_partial_sum22(reg_psum12_23_2), .reg_weight21(reg_weight12_23_1), .reg_weight22(reg_weight12_23_2), .reg_activation12(reg_activation12_23_1), .reg_activation22(reg_activation12_23_2), .weight_en(weight_en));
SA22 U12_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_24_1), .partial_sum_in12(reg_psum11_24_2), .weight_in11(reg_weight11_24_1), .weight_in12(reg_weight11_24_2), .activation_in11(reg_activation12_23_1), .activation_in21(reg_activation12_23_2), .reg_partial_sum21(reg_psum12_24_1), .reg_partial_sum22(reg_psum12_24_2), .reg_weight21(reg_weight12_24_1), .reg_weight22(reg_weight12_24_2), .reg_activation12(reg_activation12_24_1), .reg_activation22(reg_activation12_24_2), .weight_en(weight_en));
SA22 U12_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_25_1), .partial_sum_in12(reg_psum11_25_2), .weight_in11(reg_weight11_25_1), .weight_in12(reg_weight11_25_2), .activation_in11(reg_activation12_24_1), .activation_in21(reg_activation12_24_2), .reg_partial_sum21(reg_psum12_25_1), .reg_partial_sum22(reg_psum12_25_2), .reg_weight21(reg_weight12_25_1), .reg_weight22(reg_weight12_25_2), .reg_activation12(reg_activation12_25_1), .reg_activation22(reg_activation12_25_2), .weight_en(weight_en));
SA22 U12_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_26_1), .partial_sum_in12(reg_psum11_26_2), .weight_in11(reg_weight11_26_1), .weight_in12(reg_weight11_26_2), .activation_in11(reg_activation12_25_1), .activation_in21(reg_activation12_25_2), .reg_partial_sum21(reg_psum12_26_1), .reg_partial_sum22(reg_psum12_26_2), .reg_weight21(reg_weight12_26_1), .reg_weight22(reg_weight12_26_2), .reg_activation12(reg_activation12_26_1), .reg_activation22(reg_activation12_26_2), .weight_en(weight_en));
SA22 U12_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_27_1), .partial_sum_in12(reg_psum11_27_2), .weight_in11(reg_weight11_27_1), .weight_in12(reg_weight11_27_2), .activation_in11(reg_activation12_26_1), .activation_in21(reg_activation12_26_2), .reg_partial_sum21(reg_psum12_27_1), .reg_partial_sum22(reg_psum12_27_2), .reg_weight21(reg_weight12_27_1), .reg_weight22(reg_weight12_27_2), .reg_activation12(reg_activation12_27_1), .reg_activation22(reg_activation12_27_2), .weight_en(weight_en));
SA22 U12_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_28_1), .partial_sum_in12(reg_psum11_28_2), .weight_in11(reg_weight11_28_1), .weight_in12(reg_weight11_28_2), .activation_in11(reg_activation12_27_1), .activation_in21(reg_activation12_27_2), .reg_partial_sum21(reg_psum12_28_1), .reg_partial_sum22(reg_psum12_28_2), .reg_weight21(reg_weight12_28_1), .reg_weight22(reg_weight12_28_2), .reg_activation12(reg_activation12_28_1), .reg_activation22(reg_activation12_28_2), .weight_en(weight_en));
SA22 U12_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_29_1), .partial_sum_in12(reg_psum11_29_2), .weight_in11(reg_weight11_29_1), .weight_in12(reg_weight11_29_2), .activation_in11(reg_activation12_28_1), .activation_in21(reg_activation12_28_2), .reg_partial_sum21(reg_psum12_29_1), .reg_partial_sum22(reg_psum12_29_2), .reg_weight21(reg_weight12_29_1), .reg_weight22(reg_weight12_29_2), .reg_activation12(reg_activation12_29_1), .reg_activation22(reg_activation12_29_2), .weight_en(weight_en));
SA22 U12_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_30_1), .partial_sum_in12(reg_psum11_30_2), .weight_in11(reg_weight11_30_1), .weight_in12(reg_weight11_30_2), .activation_in11(reg_activation12_29_1), .activation_in21(reg_activation12_29_2), .reg_partial_sum21(reg_psum12_30_1), .reg_partial_sum22(reg_psum12_30_2), .reg_weight21(reg_weight12_30_1), .reg_weight22(reg_weight12_30_2), .reg_activation12(reg_activation12_30_1), .reg_activation22(reg_activation12_30_2), .weight_en(weight_en));
SA22 U12_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_31_1), .partial_sum_in12(reg_psum11_31_2), .weight_in11(reg_weight11_31_1), .weight_in12(reg_weight11_31_2), .activation_in11(reg_activation12_30_1), .activation_in21(reg_activation12_30_2), .reg_partial_sum21(reg_psum12_31_1), .reg_partial_sum22(reg_psum12_31_2), .reg_weight21(reg_weight12_31_1), .reg_weight22(reg_weight12_31_2), .reg_activation12(reg_activation12_31_1), .reg_activation22(reg_activation12_31_2), .weight_en(weight_en));
SA22 U12_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum11_32_1), .partial_sum_in12(reg_psum11_32_2), .weight_in11(reg_weight11_32_1), .weight_in12(reg_weight11_32_2), .activation_in11(reg_activation12_31_1), .activation_in21(reg_activation12_31_2), .reg_partial_sum21(reg_psum12_32_1), .reg_partial_sum22(reg_psum12_32_2), .reg_weight21(reg_weight12_32_1), .reg_weight22(reg_weight12_32_2), .weight_en(weight_en));
SA22 U13_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_1_1), .partial_sum_in12(reg_psum12_1_2), .weight_in11(reg_weight12_1_1), .weight_in12(reg_weight12_1_2), .activation_in11(in_activation13_1_1), .activation_in21(in_activation13_1_2), .reg_partial_sum21(reg_psum13_1_1), .reg_partial_sum22(reg_psum13_1_2), .reg_weight21(reg_weight13_1_1), .reg_weight22(reg_weight13_1_2), .reg_activation12(reg_activation13_1_1), .reg_activation22(reg_activation13_1_2), .weight_en(weight_en));
SA22 U13_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_2_1), .partial_sum_in12(reg_psum12_2_2), .weight_in11(reg_weight12_2_1), .weight_in12(reg_weight12_2_2), .activation_in11(reg_activation13_1_1), .activation_in21(reg_activation13_1_2), .reg_partial_sum21(reg_psum13_2_1), .reg_partial_sum22(reg_psum13_2_2), .reg_weight21(reg_weight13_2_1), .reg_weight22(reg_weight13_2_2), .reg_activation12(reg_activation13_2_1), .reg_activation22(reg_activation13_2_2), .weight_en(weight_en));
SA22 U13_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_3_1), .partial_sum_in12(reg_psum12_3_2), .weight_in11(reg_weight12_3_1), .weight_in12(reg_weight12_3_2), .activation_in11(reg_activation13_2_1), .activation_in21(reg_activation13_2_2), .reg_partial_sum21(reg_psum13_3_1), .reg_partial_sum22(reg_psum13_3_2), .reg_weight21(reg_weight13_3_1), .reg_weight22(reg_weight13_3_2), .reg_activation12(reg_activation13_3_1), .reg_activation22(reg_activation13_3_2), .weight_en(weight_en));
SA22 U13_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_4_1), .partial_sum_in12(reg_psum12_4_2), .weight_in11(reg_weight12_4_1), .weight_in12(reg_weight12_4_2), .activation_in11(reg_activation13_3_1), .activation_in21(reg_activation13_3_2), .reg_partial_sum21(reg_psum13_4_1), .reg_partial_sum22(reg_psum13_4_2), .reg_weight21(reg_weight13_4_1), .reg_weight22(reg_weight13_4_2), .reg_activation12(reg_activation13_4_1), .reg_activation22(reg_activation13_4_2), .weight_en(weight_en));
SA22 U13_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_5_1), .partial_sum_in12(reg_psum12_5_2), .weight_in11(reg_weight12_5_1), .weight_in12(reg_weight12_5_2), .activation_in11(reg_activation13_4_1), .activation_in21(reg_activation13_4_2), .reg_partial_sum21(reg_psum13_5_1), .reg_partial_sum22(reg_psum13_5_2), .reg_weight21(reg_weight13_5_1), .reg_weight22(reg_weight13_5_2), .reg_activation12(reg_activation13_5_1), .reg_activation22(reg_activation13_5_2), .weight_en(weight_en));
SA22 U13_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_6_1), .partial_sum_in12(reg_psum12_6_2), .weight_in11(reg_weight12_6_1), .weight_in12(reg_weight12_6_2), .activation_in11(reg_activation13_5_1), .activation_in21(reg_activation13_5_2), .reg_partial_sum21(reg_psum13_6_1), .reg_partial_sum22(reg_psum13_6_2), .reg_weight21(reg_weight13_6_1), .reg_weight22(reg_weight13_6_2), .reg_activation12(reg_activation13_6_1), .reg_activation22(reg_activation13_6_2), .weight_en(weight_en));
SA22 U13_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_7_1), .partial_sum_in12(reg_psum12_7_2), .weight_in11(reg_weight12_7_1), .weight_in12(reg_weight12_7_2), .activation_in11(reg_activation13_6_1), .activation_in21(reg_activation13_6_2), .reg_partial_sum21(reg_psum13_7_1), .reg_partial_sum22(reg_psum13_7_2), .reg_weight21(reg_weight13_7_1), .reg_weight22(reg_weight13_7_2), .reg_activation12(reg_activation13_7_1), .reg_activation22(reg_activation13_7_2), .weight_en(weight_en));
SA22 U13_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_8_1), .partial_sum_in12(reg_psum12_8_2), .weight_in11(reg_weight12_8_1), .weight_in12(reg_weight12_8_2), .activation_in11(reg_activation13_7_1), .activation_in21(reg_activation13_7_2), .reg_partial_sum21(reg_psum13_8_1), .reg_partial_sum22(reg_psum13_8_2), .reg_weight21(reg_weight13_8_1), .reg_weight22(reg_weight13_8_2), .reg_activation12(reg_activation13_8_1), .reg_activation22(reg_activation13_8_2), .weight_en(weight_en));
SA22 U13_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_9_1), .partial_sum_in12(reg_psum12_9_2), .weight_in11(reg_weight12_9_1), .weight_in12(reg_weight12_9_2), .activation_in11(reg_activation13_8_1), .activation_in21(reg_activation13_8_2), .reg_partial_sum21(reg_psum13_9_1), .reg_partial_sum22(reg_psum13_9_2), .reg_weight21(reg_weight13_9_1), .reg_weight22(reg_weight13_9_2), .reg_activation12(reg_activation13_9_1), .reg_activation22(reg_activation13_9_2), .weight_en(weight_en));
SA22 U13_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_10_1), .partial_sum_in12(reg_psum12_10_2), .weight_in11(reg_weight12_10_1), .weight_in12(reg_weight12_10_2), .activation_in11(reg_activation13_9_1), .activation_in21(reg_activation13_9_2), .reg_partial_sum21(reg_psum13_10_1), .reg_partial_sum22(reg_psum13_10_2), .reg_weight21(reg_weight13_10_1), .reg_weight22(reg_weight13_10_2), .reg_activation12(reg_activation13_10_1), .reg_activation22(reg_activation13_10_2), .weight_en(weight_en));
SA22 U13_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_11_1), .partial_sum_in12(reg_psum12_11_2), .weight_in11(reg_weight12_11_1), .weight_in12(reg_weight12_11_2), .activation_in11(reg_activation13_10_1), .activation_in21(reg_activation13_10_2), .reg_partial_sum21(reg_psum13_11_1), .reg_partial_sum22(reg_psum13_11_2), .reg_weight21(reg_weight13_11_1), .reg_weight22(reg_weight13_11_2), .reg_activation12(reg_activation13_11_1), .reg_activation22(reg_activation13_11_2), .weight_en(weight_en));
SA22 U13_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_12_1), .partial_sum_in12(reg_psum12_12_2), .weight_in11(reg_weight12_12_1), .weight_in12(reg_weight12_12_2), .activation_in11(reg_activation13_11_1), .activation_in21(reg_activation13_11_2), .reg_partial_sum21(reg_psum13_12_1), .reg_partial_sum22(reg_psum13_12_2), .reg_weight21(reg_weight13_12_1), .reg_weight22(reg_weight13_12_2), .reg_activation12(reg_activation13_12_1), .reg_activation22(reg_activation13_12_2), .weight_en(weight_en));
SA22 U13_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_13_1), .partial_sum_in12(reg_psum12_13_2), .weight_in11(reg_weight12_13_1), .weight_in12(reg_weight12_13_2), .activation_in11(reg_activation13_12_1), .activation_in21(reg_activation13_12_2), .reg_partial_sum21(reg_psum13_13_1), .reg_partial_sum22(reg_psum13_13_2), .reg_weight21(reg_weight13_13_1), .reg_weight22(reg_weight13_13_2), .reg_activation12(reg_activation13_13_1), .reg_activation22(reg_activation13_13_2), .weight_en(weight_en));
SA22 U13_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_14_1), .partial_sum_in12(reg_psum12_14_2), .weight_in11(reg_weight12_14_1), .weight_in12(reg_weight12_14_2), .activation_in11(reg_activation13_13_1), .activation_in21(reg_activation13_13_2), .reg_partial_sum21(reg_psum13_14_1), .reg_partial_sum22(reg_psum13_14_2), .reg_weight21(reg_weight13_14_1), .reg_weight22(reg_weight13_14_2), .reg_activation12(reg_activation13_14_1), .reg_activation22(reg_activation13_14_2), .weight_en(weight_en));
SA22 U13_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_15_1), .partial_sum_in12(reg_psum12_15_2), .weight_in11(reg_weight12_15_1), .weight_in12(reg_weight12_15_2), .activation_in11(reg_activation13_14_1), .activation_in21(reg_activation13_14_2), .reg_partial_sum21(reg_psum13_15_1), .reg_partial_sum22(reg_psum13_15_2), .reg_weight21(reg_weight13_15_1), .reg_weight22(reg_weight13_15_2), .reg_activation12(reg_activation13_15_1), .reg_activation22(reg_activation13_15_2), .weight_en(weight_en));
SA22 U13_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_16_1), .partial_sum_in12(reg_psum12_16_2), .weight_in11(reg_weight12_16_1), .weight_in12(reg_weight12_16_2), .activation_in11(reg_activation13_15_1), .activation_in21(reg_activation13_15_2), .reg_partial_sum21(reg_psum13_16_1), .reg_partial_sum22(reg_psum13_16_2), .reg_weight21(reg_weight13_16_1), .reg_weight22(reg_weight13_16_2), .reg_activation12(reg_activation13_16_1), .reg_activation22(reg_activation13_16_2), .weight_en(weight_en));
SA22 U13_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_17_1), .partial_sum_in12(reg_psum12_17_2), .weight_in11(reg_weight12_17_1), .weight_in12(reg_weight12_17_2), .activation_in11(reg_activation13_16_1), .activation_in21(reg_activation13_16_2), .reg_partial_sum21(reg_psum13_17_1), .reg_partial_sum22(reg_psum13_17_2), .reg_weight21(reg_weight13_17_1), .reg_weight22(reg_weight13_17_2), .reg_activation12(reg_activation13_17_1), .reg_activation22(reg_activation13_17_2), .weight_en(weight_en));
SA22 U13_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_18_1), .partial_sum_in12(reg_psum12_18_2), .weight_in11(reg_weight12_18_1), .weight_in12(reg_weight12_18_2), .activation_in11(reg_activation13_17_1), .activation_in21(reg_activation13_17_2), .reg_partial_sum21(reg_psum13_18_1), .reg_partial_sum22(reg_psum13_18_2), .reg_weight21(reg_weight13_18_1), .reg_weight22(reg_weight13_18_2), .reg_activation12(reg_activation13_18_1), .reg_activation22(reg_activation13_18_2), .weight_en(weight_en));
SA22 U13_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_19_1), .partial_sum_in12(reg_psum12_19_2), .weight_in11(reg_weight12_19_1), .weight_in12(reg_weight12_19_2), .activation_in11(reg_activation13_18_1), .activation_in21(reg_activation13_18_2), .reg_partial_sum21(reg_psum13_19_1), .reg_partial_sum22(reg_psum13_19_2), .reg_weight21(reg_weight13_19_1), .reg_weight22(reg_weight13_19_2), .reg_activation12(reg_activation13_19_1), .reg_activation22(reg_activation13_19_2), .weight_en(weight_en));
SA22 U13_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_20_1), .partial_sum_in12(reg_psum12_20_2), .weight_in11(reg_weight12_20_1), .weight_in12(reg_weight12_20_2), .activation_in11(reg_activation13_19_1), .activation_in21(reg_activation13_19_2), .reg_partial_sum21(reg_psum13_20_1), .reg_partial_sum22(reg_psum13_20_2), .reg_weight21(reg_weight13_20_1), .reg_weight22(reg_weight13_20_2), .reg_activation12(reg_activation13_20_1), .reg_activation22(reg_activation13_20_2), .weight_en(weight_en));
SA22 U13_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_21_1), .partial_sum_in12(reg_psum12_21_2), .weight_in11(reg_weight12_21_1), .weight_in12(reg_weight12_21_2), .activation_in11(reg_activation13_20_1), .activation_in21(reg_activation13_20_2), .reg_partial_sum21(reg_psum13_21_1), .reg_partial_sum22(reg_psum13_21_2), .reg_weight21(reg_weight13_21_1), .reg_weight22(reg_weight13_21_2), .reg_activation12(reg_activation13_21_1), .reg_activation22(reg_activation13_21_2), .weight_en(weight_en));
SA22 U13_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_22_1), .partial_sum_in12(reg_psum12_22_2), .weight_in11(reg_weight12_22_1), .weight_in12(reg_weight12_22_2), .activation_in11(reg_activation13_21_1), .activation_in21(reg_activation13_21_2), .reg_partial_sum21(reg_psum13_22_1), .reg_partial_sum22(reg_psum13_22_2), .reg_weight21(reg_weight13_22_1), .reg_weight22(reg_weight13_22_2), .reg_activation12(reg_activation13_22_1), .reg_activation22(reg_activation13_22_2), .weight_en(weight_en));
SA22 U13_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_23_1), .partial_sum_in12(reg_psum12_23_2), .weight_in11(reg_weight12_23_1), .weight_in12(reg_weight12_23_2), .activation_in11(reg_activation13_22_1), .activation_in21(reg_activation13_22_2), .reg_partial_sum21(reg_psum13_23_1), .reg_partial_sum22(reg_psum13_23_2), .reg_weight21(reg_weight13_23_1), .reg_weight22(reg_weight13_23_2), .reg_activation12(reg_activation13_23_1), .reg_activation22(reg_activation13_23_2), .weight_en(weight_en));
SA22 U13_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_24_1), .partial_sum_in12(reg_psum12_24_2), .weight_in11(reg_weight12_24_1), .weight_in12(reg_weight12_24_2), .activation_in11(reg_activation13_23_1), .activation_in21(reg_activation13_23_2), .reg_partial_sum21(reg_psum13_24_1), .reg_partial_sum22(reg_psum13_24_2), .reg_weight21(reg_weight13_24_1), .reg_weight22(reg_weight13_24_2), .reg_activation12(reg_activation13_24_1), .reg_activation22(reg_activation13_24_2), .weight_en(weight_en));
SA22 U13_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_25_1), .partial_sum_in12(reg_psum12_25_2), .weight_in11(reg_weight12_25_1), .weight_in12(reg_weight12_25_2), .activation_in11(reg_activation13_24_1), .activation_in21(reg_activation13_24_2), .reg_partial_sum21(reg_psum13_25_1), .reg_partial_sum22(reg_psum13_25_2), .reg_weight21(reg_weight13_25_1), .reg_weight22(reg_weight13_25_2), .reg_activation12(reg_activation13_25_1), .reg_activation22(reg_activation13_25_2), .weight_en(weight_en));
SA22 U13_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_26_1), .partial_sum_in12(reg_psum12_26_2), .weight_in11(reg_weight12_26_1), .weight_in12(reg_weight12_26_2), .activation_in11(reg_activation13_25_1), .activation_in21(reg_activation13_25_2), .reg_partial_sum21(reg_psum13_26_1), .reg_partial_sum22(reg_psum13_26_2), .reg_weight21(reg_weight13_26_1), .reg_weight22(reg_weight13_26_2), .reg_activation12(reg_activation13_26_1), .reg_activation22(reg_activation13_26_2), .weight_en(weight_en));
SA22 U13_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_27_1), .partial_sum_in12(reg_psum12_27_2), .weight_in11(reg_weight12_27_1), .weight_in12(reg_weight12_27_2), .activation_in11(reg_activation13_26_1), .activation_in21(reg_activation13_26_2), .reg_partial_sum21(reg_psum13_27_1), .reg_partial_sum22(reg_psum13_27_2), .reg_weight21(reg_weight13_27_1), .reg_weight22(reg_weight13_27_2), .reg_activation12(reg_activation13_27_1), .reg_activation22(reg_activation13_27_2), .weight_en(weight_en));
SA22 U13_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_28_1), .partial_sum_in12(reg_psum12_28_2), .weight_in11(reg_weight12_28_1), .weight_in12(reg_weight12_28_2), .activation_in11(reg_activation13_27_1), .activation_in21(reg_activation13_27_2), .reg_partial_sum21(reg_psum13_28_1), .reg_partial_sum22(reg_psum13_28_2), .reg_weight21(reg_weight13_28_1), .reg_weight22(reg_weight13_28_2), .reg_activation12(reg_activation13_28_1), .reg_activation22(reg_activation13_28_2), .weight_en(weight_en));
SA22 U13_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_29_1), .partial_sum_in12(reg_psum12_29_2), .weight_in11(reg_weight12_29_1), .weight_in12(reg_weight12_29_2), .activation_in11(reg_activation13_28_1), .activation_in21(reg_activation13_28_2), .reg_partial_sum21(reg_psum13_29_1), .reg_partial_sum22(reg_psum13_29_2), .reg_weight21(reg_weight13_29_1), .reg_weight22(reg_weight13_29_2), .reg_activation12(reg_activation13_29_1), .reg_activation22(reg_activation13_29_2), .weight_en(weight_en));
SA22 U13_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_30_1), .partial_sum_in12(reg_psum12_30_2), .weight_in11(reg_weight12_30_1), .weight_in12(reg_weight12_30_2), .activation_in11(reg_activation13_29_1), .activation_in21(reg_activation13_29_2), .reg_partial_sum21(reg_psum13_30_1), .reg_partial_sum22(reg_psum13_30_2), .reg_weight21(reg_weight13_30_1), .reg_weight22(reg_weight13_30_2), .reg_activation12(reg_activation13_30_1), .reg_activation22(reg_activation13_30_2), .weight_en(weight_en));
SA22 U13_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_31_1), .partial_sum_in12(reg_psum12_31_2), .weight_in11(reg_weight12_31_1), .weight_in12(reg_weight12_31_2), .activation_in11(reg_activation13_30_1), .activation_in21(reg_activation13_30_2), .reg_partial_sum21(reg_psum13_31_1), .reg_partial_sum22(reg_psum13_31_2), .reg_weight21(reg_weight13_31_1), .reg_weight22(reg_weight13_31_2), .reg_activation12(reg_activation13_31_1), .reg_activation22(reg_activation13_31_2), .weight_en(weight_en));
SA22 U13_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum12_32_1), .partial_sum_in12(reg_psum12_32_2), .weight_in11(reg_weight12_32_1), .weight_in12(reg_weight12_32_2), .activation_in11(reg_activation13_31_1), .activation_in21(reg_activation13_31_2), .reg_partial_sum21(reg_psum13_32_1), .reg_partial_sum22(reg_psum13_32_2), .reg_weight21(reg_weight13_32_1), .reg_weight22(reg_weight13_32_2), .weight_en(weight_en));
SA22 U14_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_1_1), .partial_sum_in12(reg_psum13_1_2), .weight_in11(reg_weight13_1_1), .weight_in12(reg_weight13_1_2), .activation_in11(in_activation14_1_1), .activation_in21(in_activation14_1_2), .reg_partial_sum21(reg_psum14_1_1), .reg_partial_sum22(reg_psum14_1_2), .reg_weight21(reg_weight14_1_1), .reg_weight22(reg_weight14_1_2), .reg_activation12(reg_activation14_1_1), .reg_activation22(reg_activation14_1_2), .weight_en(weight_en));
SA22 U14_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_2_1), .partial_sum_in12(reg_psum13_2_2), .weight_in11(reg_weight13_2_1), .weight_in12(reg_weight13_2_2), .activation_in11(reg_activation14_1_1), .activation_in21(reg_activation14_1_2), .reg_partial_sum21(reg_psum14_2_1), .reg_partial_sum22(reg_psum14_2_2), .reg_weight21(reg_weight14_2_1), .reg_weight22(reg_weight14_2_2), .reg_activation12(reg_activation14_2_1), .reg_activation22(reg_activation14_2_2), .weight_en(weight_en));
SA22 U14_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_3_1), .partial_sum_in12(reg_psum13_3_2), .weight_in11(reg_weight13_3_1), .weight_in12(reg_weight13_3_2), .activation_in11(reg_activation14_2_1), .activation_in21(reg_activation14_2_2), .reg_partial_sum21(reg_psum14_3_1), .reg_partial_sum22(reg_psum14_3_2), .reg_weight21(reg_weight14_3_1), .reg_weight22(reg_weight14_3_2), .reg_activation12(reg_activation14_3_1), .reg_activation22(reg_activation14_3_2), .weight_en(weight_en));
SA22 U14_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_4_1), .partial_sum_in12(reg_psum13_4_2), .weight_in11(reg_weight13_4_1), .weight_in12(reg_weight13_4_2), .activation_in11(reg_activation14_3_1), .activation_in21(reg_activation14_3_2), .reg_partial_sum21(reg_psum14_4_1), .reg_partial_sum22(reg_psum14_4_2), .reg_weight21(reg_weight14_4_1), .reg_weight22(reg_weight14_4_2), .reg_activation12(reg_activation14_4_1), .reg_activation22(reg_activation14_4_2), .weight_en(weight_en));
SA22 U14_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_5_1), .partial_sum_in12(reg_psum13_5_2), .weight_in11(reg_weight13_5_1), .weight_in12(reg_weight13_5_2), .activation_in11(reg_activation14_4_1), .activation_in21(reg_activation14_4_2), .reg_partial_sum21(reg_psum14_5_1), .reg_partial_sum22(reg_psum14_5_2), .reg_weight21(reg_weight14_5_1), .reg_weight22(reg_weight14_5_2), .reg_activation12(reg_activation14_5_1), .reg_activation22(reg_activation14_5_2), .weight_en(weight_en));
SA22 U14_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_6_1), .partial_sum_in12(reg_psum13_6_2), .weight_in11(reg_weight13_6_1), .weight_in12(reg_weight13_6_2), .activation_in11(reg_activation14_5_1), .activation_in21(reg_activation14_5_2), .reg_partial_sum21(reg_psum14_6_1), .reg_partial_sum22(reg_psum14_6_2), .reg_weight21(reg_weight14_6_1), .reg_weight22(reg_weight14_6_2), .reg_activation12(reg_activation14_6_1), .reg_activation22(reg_activation14_6_2), .weight_en(weight_en));
SA22 U14_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_7_1), .partial_sum_in12(reg_psum13_7_2), .weight_in11(reg_weight13_7_1), .weight_in12(reg_weight13_7_2), .activation_in11(reg_activation14_6_1), .activation_in21(reg_activation14_6_2), .reg_partial_sum21(reg_psum14_7_1), .reg_partial_sum22(reg_psum14_7_2), .reg_weight21(reg_weight14_7_1), .reg_weight22(reg_weight14_7_2), .reg_activation12(reg_activation14_7_1), .reg_activation22(reg_activation14_7_2), .weight_en(weight_en));
SA22 U14_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_8_1), .partial_sum_in12(reg_psum13_8_2), .weight_in11(reg_weight13_8_1), .weight_in12(reg_weight13_8_2), .activation_in11(reg_activation14_7_1), .activation_in21(reg_activation14_7_2), .reg_partial_sum21(reg_psum14_8_1), .reg_partial_sum22(reg_psum14_8_2), .reg_weight21(reg_weight14_8_1), .reg_weight22(reg_weight14_8_2), .reg_activation12(reg_activation14_8_1), .reg_activation22(reg_activation14_8_2), .weight_en(weight_en));
SA22 U14_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_9_1), .partial_sum_in12(reg_psum13_9_2), .weight_in11(reg_weight13_9_1), .weight_in12(reg_weight13_9_2), .activation_in11(reg_activation14_8_1), .activation_in21(reg_activation14_8_2), .reg_partial_sum21(reg_psum14_9_1), .reg_partial_sum22(reg_psum14_9_2), .reg_weight21(reg_weight14_9_1), .reg_weight22(reg_weight14_9_2), .reg_activation12(reg_activation14_9_1), .reg_activation22(reg_activation14_9_2), .weight_en(weight_en));
SA22 U14_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_10_1), .partial_sum_in12(reg_psum13_10_2), .weight_in11(reg_weight13_10_1), .weight_in12(reg_weight13_10_2), .activation_in11(reg_activation14_9_1), .activation_in21(reg_activation14_9_2), .reg_partial_sum21(reg_psum14_10_1), .reg_partial_sum22(reg_psum14_10_2), .reg_weight21(reg_weight14_10_1), .reg_weight22(reg_weight14_10_2), .reg_activation12(reg_activation14_10_1), .reg_activation22(reg_activation14_10_2), .weight_en(weight_en));
SA22 U14_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_11_1), .partial_sum_in12(reg_psum13_11_2), .weight_in11(reg_weight13_11_1), .weight_in12(reg_weight13_11_2), .activation_in11(reg_activation14_10_1), .activation_in21(reg_activation14_10_2), .reg_partial_sum21(reg_psum14_11_1), .reg_partial_sum22(reg_psum14_11_2), .reg_weight21(reg_weight14_11_1), .reg_weight22(reg_weight14_11_2), .reg_activation12(reg_activation14_11_1), .reg_activation22(reg_activation14_11_2), .weight_en(weight_en));
SA22 U14_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_12_1), .partial_sum_in12(reg_psum13_12_2), .weight_in11(reg_weight13_12_1), .weight_in12(reg_weight13_12_2), .activation_in11(reg_activation14_11_1), .activation_in21(reg_activation14_11_2), .reg_partial_sum21(reg_psum14_12_1), .reg_partial_sum22(reg_psum14_12_2), .reg_weight21(reg_weight14_12_1), .reg_weight22(reg_weight14_12_2), .reg_activation12(reg_activation14_12_1), .reg_activation22(reg_activation14_12_2), .weight_en(weight_en));
SA22 U14_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_13_1), .partial_sum_in12(reg_psum13_13_2), .weight_in11(reg_weight13_13_1), .weight_in12(reg_weight13_13_2), .activation_in11(reg_activation14_12_1), .activation_in21(reg_activation14_12_2), .reg_partial_sum21(reg_psum14_13_1), .reg_partial_sum22(reg_psum14_13_2), .reg_weight21(reg_weight14_13_1), .reg_weight22(reg_weight14_13_2), .reg_activation12(reg_activation14_13_1), .reg_activation22(reg_activation14_13_2), .weight_en(weight_en));
SA22 U14_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_14_1), .partial_sum_in12(reg_psum13_14_2), .weight_in11(reg_weight13_14_1), .weight_in12(reg_weight13_14_2), .activation_in11(reg_activation14_13_1), .activation_in21(reg_activation14_13_2), .reg_partial_sum21(reg_psum14_14_1), .reg_partial_sum22(reg_psum14_14_2), .reg_weight21(reg_weight14_14_1), .reg_weight22(reg_weight14_14_2), .reg_activation12(reg_activation14_14_1), .reg_activation22(reg_activation14_14_2), .weight_en(weight_en));
SA22 U14_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_15_1), .partial_sum_in12(reg_psum13_15_2), .weight_in11(reg_weight13_15_1), .weight_in12(reg_weight13_15_2), .activation_in11(reg_activation14_14_1), .activation_in21(reg_activation14_14_2), .reg_partial_sum21(reg_psum14_15_1), .reg_partial_sum22(reg_psum14_15_2), .reg_weight21(reg_weight14_15_1), .reg_weight22(reg_weight14_15_2), .reg_activation12(reg_activation14_15_1), .reg_activation22(reg_activation14_15_2), .weight_en(weight_en));
SA22 U14_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_16_1), .partial_sum_in12(reg_psum13_16_2), .weight_in11(reg_weight13_16_1), .weight_in12(reg_weight13_16_2), .activation_in11(reg_activation14_15_1), .activation_in21(reg_activation14_15_2), .reg_partial_sum21(reg_psum14_16_1), .reg_partial_sum22(reg_psum14_16_2), .reg_weight21(reg_weight14_16_1), .reg_weight22(reg_weight14_16_2), .reg_activation12(reg_activation14_16_1), .reg_activation22(reg_activation14_16_2), .weight_en(weight_en));
SA22 U14_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_17_1), .partial_sum_in12(reg_psum13_17_2), .weight_in11(reg_weight13_17_1), .weight_in12(reg_weight13_17_2), .activation_in11(reg_activation14_16_1), .activation_in21(reg_activation14_16_2), .reg_partial_sum21(reg_psum14_17_1), .reg_partial_sum22(reg_psum14_17_2), .reg_weight21(reg_weight14_17_1), .reg_weight22(reg_weight14_17_2), .reg_activation12(reg_activation14_17_1), .reg_activation22(reg_activation14_17_2), .weight_en(weight_en));
SA22 U14_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_18_1), .partial_sum_in12(reg_psum13_18_2), .weight_in11(reg_weight13_18_1), .weight_in12(reg_weight13_18_2), .activation_in11(reg_activation14_17_1), .activation_in21(reg_activation14_17_2), .reg_partial_sum21(reg_psum14_18_1), .reg_partial_sum22(reg_psum14_18_2), .reg_weight21(reg_weight14_18_1), .reg_weight22(reg_weight14_18_2), .reg_activation12(reg_activation14_18_1), .reg_activation22(reg_activation14_18_2), .weight_en(weight_en));
SA22 U14_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_19_1), .partial_sum_in12(reg_psum13_19_2), .weight_in11(reg_weight13_19_1), .weight_in12(reg_weight13_19_2), .activation_in11(reg_activation14_18_1), .activation_in21(reg_activation14_18_2), .reg_partial_sum21(reg_psum14_19_1), .reg_partial_sum22(reg_psum14_19_2), .reg_weight21(reg_weight14_19_1), .reg_weight22(reg_weight14_19_2), .reg_activation12(reg_activation14_19_1), .reg_activation22(reg_activation14_19_2), .weight_en(weight_en));
SA22 U14_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_20_1), .partial_sum_in12(reg_psum13_20_2), .weight_in11(reg_weight13_20_1), .weight_in12(reg_weight13_20_2), .activation_in11(reg_activation14_19_1), .activation_in21(reg_activation14_19_2), .reg_partial_sum21(reg_psum14_20_1), .reg_partial_sum22(reg_psum14_20_2), .reg_weight21(reg_weight14_20_1), .reg_weight22(reg_weight14_20_2), .reg_activation12(reg_activation14_20_1), .reg_activation22(reg_activation14_20_2), .weight_en(weight_en));
SA22 U14_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_21_1), .partial_sum_in12(reg_psum13_21_2), .weight_in11(reg_weight13_21_1), .weight_in12(reg_weight13_21_2), .activation_in11(reg_activation14_20_1), .activation_in21(reg_activation14_20_2), .reg_partial_sum21(reg_psum14_21_1), .reg_partial_sum22(reg_psum14_21_2), .reg_weight21(reg_weight14_21_1), .reg_weight22(reg_weight14_21_2), .reg_activation12(reg_activation14_21_1), .reg_activation22(reg_activation14_21_2), .weight_en(weight_en));
SA22 U14_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_22_1), .partial_sum_in12(reg_psum13_22_2), .weight_in11(reg_weight13_22_1), .weight_in12(reg_weight13_22_2), .activation_in11(reg_activation14_21_1), .activation_in21(reg_activation14_21_2), .reg_partial_sum21(reg_psum14_22_1), .reg_partial_sum22(reg_psum14_22_2), .reg_weight21(reg_weight14_22_1), .reg_weight22(reg_weight14_22_2), .reg_activation12(reg_activation14_22_1), .reg_activation22(reg_activation14_22_2), .weight_en(weight_en));
SA22 U14_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_23_1), .partial_sum_in12(reg_psum13_23_2), .weight_in11(reg_weight13_23_1), .weight_in12(reg_weight13_23_2), .activation_in11(reg_activation14_22_1), .activation_in21(reg_activation14_22_2), .reg_partial_sum21(reg_psum14_23_1), .reg_partial_sum22(reg_psum14_23_2), .reg_weight21(reg_weight14_23_1), .reg_weight22(reg_weight14_23_2), .reg_activation12(reg_activation14_23_1), .reg_activation22(reg_activation14_23_2), .weight_en(weight_en));
SA22 U14_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_24_1), .partial_sum_in12(reg_psum13_24_2), .weight_in11(reg_weight13_24_1), .weight_in12(reg_weight13_24_2), .activation_in11(reg_activation14_23_1), .activation_in21(reg_activation14_23_2), .reg_partial_sum21(reg_psum14_24_1), .reg_partial_sum22(reg_psum14_24_2), .reg_weight21(reg_weight14_24_1), .reg_weight22(reg_weight14_24_2), .reg_activation12(reg_activation14_24_1), .reg_activation22(reg_activation14_24_2), .weight_en(weight_en));
SA22 U14_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_25_1), .partial_sum_in12(reg_psum13_25_2), .weight_in11(reg_weight13_25_1), .weight_in12(reg_weight13_25_2), .activation_in11(reg_activation14_24_1), .activation_in21(reg_activation14_24_2), .reg_partial_sum21(reg_psum14_25_1), .reg_partial_sum22(reg_psum14_25_2), .reg_weight21(reg_weight14_25_1), .reg_weight22(reg_weight14_25_2), .reg_activation12(reg_activation14_25_1), .reg_activation22(reg_activation14_25_2), .weight_en(weight_en));
SA22 U14_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_26_1), .partial_sum_in12(reg_psum13_26_2), .weight_in11(reg_weight13_26_1), .weight_in12(reg_weight13_26_2), .activation_in11(reg_activation14_25_1), .activation_in21(reg_activation14_25_2), .reg_partial_sum21(reg_psum14_26_1), .reg_partial_sum22(reg_psum14_26_2), .reg_weight21(reg_weight14_26_1), .reg_weight22(reg_weight14_26_2), .reg_activation12(reg_activation14_26_1), .reg_activation22(reg_activation14_26_2), .weight_en(weight_en));
SA22 U14_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_27_1), .partial_sum_in12(reg_psum13_27_2), .weight_in11(reg_weight13_27_1), .weight_in12(reg_weight13_27_2), .activation_in11(reg_activation14_26_1), .activation_in21(reg_activation14_26_2), .reg_partial_sum21(reg_psum14_27_1), .reg_partial_sum22(reg_psum14_27_2), .reg_weight21(reg_weight14_27_1), .reg_weight22(reg_weight14_27_2), .reg_activation12(reg_activation14_27_1), .reg_activation22(reg_activation14_27_2), .weight_en(weight_en));
SA22 U14_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_28_1), .partial_sum_in12(reg_psum13_28_2), .weight_in11(reg_weight13_28_1), .weight_in12(reg_weight13_28_2), .activation_in11(reg_activation14_27_1), .activation_in21(reg_activation14_27_2), .reg_partial_sum21(reg_psum14_28_1), .reg_partial_sum22(reg_psum14_28_2), .reg_weight21(reg_weight14_28_1), .reg_weight22(reg_weight14_28_2), .reg_activation12(reg_activation14_28_1), .reg_activation22(reg_activation14_28_2), .weight_en(weight_en));
SA22 U14_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_29_1), .partial_sum_in12(reg_psum13_29_2), .weight_in11(reg_weight13_29_1), .weight_in12(reg_weight13_29_2), .activation_in11(reg_activation14_28_1), .activation_in21(reg_activation14_28_2), .reg_partial_sum21(reg_psum14_29_1), .reg_partial_sum22(reg_psum14_29_2), .reg_weight21(reg_weight14_29_1), .reg_weight22(reg_weight14_29_2), .reg_activation12(reg_activation14_29_1), .reg_activation22(reg_activation14_29_2), .weight_en(weight_en));
SA22 U14_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_30_1), .partial_sum_in12(reg_psum13_30_2), .weight_in11(reg_weight13_30_1), .weight_in12(reg_weight13_30_2), .activation_in11(reg_activation14_29_1), .activation_in21(reg_activation14_29_2), .reg_partial_sum21(reg_psum14_30_1), .reg_partial_sum22(reg_psum14_30_2), .reg_weight21(reg_weight14_30_1), .reg_weight22(reg_weight14_30_2), .reg_activation12(reg_activation14_30_1), .reg_activation22(reg_activation14_30_2), .weight_en(weight_en));
SA22 U14_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_31_1), .partial_sum_in12(reg_psum13_31_2), .weight_in11(reg_weight13_31_1), .weight_in12(reg_weight13_31_2), .activation_in11(reg_activation14_30_1), .activation_in21(reg_activation14_30_2), .reg_partial_sum21(reg_psum14_31_1), .reg_partial_sum22(reg_psum14_31_2), .reg_weight21(reg_weight14_31_1), .reg_weight22(reg_weight14_31_2), .reg_activation12(reg_activation14_31_1), .reg_activation22(reg_activation14_31_2), .weight_en(weight_en));
SA22 U14_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum13_32_1), .partial_sum_in12(reg_psum13_32_2), .weight_in11(reg_weight13_32_1), .weight_in12(reg_weight13_32_2), .activation_in11(reg_activation14_31_1), .activation_in21(reg_activation14_31_2), .reg_partial_sum21(reg_psum14_32_1), .reg_partial_sum22(reg_psum14_32_2), .reg_weight21(reg_weight14_32_1), .reg_weight22(reg_weight14_32_2), .weight_en(weight_en));
SA22 U15_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_1_1), .partial_sum_in12(reg_psum14_1_2), .weight_in11(reg_weight14_1_1), .weight_in12(reg_weight14_1_2), .activation_in11(in_activation15_1_1), .activation_in21(in_activation15_1_2), .reg_partial_sum21(reg_psum15_1_1), .reg_partial_sum22(reg_psum15_1_2), .reg_weight21(reg_weight15_1_1), .reg_weight22(reg_weight15_1_2), .reg_activation12(reg_activation15_1_1), .reg_activation22(reg_activation15_1_2), .weight_en(weight_en));
SA22 U15_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_2_1), .partial_sum_in12(reg_psum14_2_2), .weight_in11(reg_weight14_2_1), .weight_in12(reg_weight14_2_2), .activation_in11(reg_activation15_1_1), .activation_in21(reg_activation15_1_2), .reg_partial_sum21(reg_psum15_2_1), .reg_partial_sum22(reg_psum15_2_2), .reg_weight21(reg_weight15_2_1), .reg_weight22(reg_weight15_2_2), .reg_activation12(reg_activation15_2_1), .reg_activation22(reg_activation15_2_2), .weight_en(weight_en));
SA22 U15_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_3_1), .partial_sum_in12(reg_psum14_3_2), .weight_in11(reg_weight14_3_1), .weight_in12(reg_weight14_3_2), .activation_in11(reg_activation15_2_1), .activation_in21(reg_activation15_2_2), .reg_partial_sum21(reg_psum15_3_1), .reg_partial_sum22(reg_psum15_3_2), .reg_weight21(reg_weight15_3_1), .reg_weight22(reg_weight15_3_2), .reg_activation12(reg_activation15_3_1), .reg_activation22(reg_activation15_3_2), .weight_en(weight_en));
SA22 U15_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_4_1), .partial_sum_in12(reg_psum14_4_2), .weight_in11(reg_weight14_4_1), .weight_in12(reg_weight14_4_2), .activation_in11(reg_activation15_3_1), .activation_in21(reg_activation15_3_2), .reg_partial_sum21(reg_psum15_4_1), .reg_partial_sum22(reg_psum15_4_2), .reg_weight21(reg_weight15_4_1), .reg_weight22(reg_weight15_4_2), .reg_activation12(reg_activation15_4_1), .reg_activation22(reg_activation15_4_2), .weight_en(weight_en));
SA22 U15_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_5_1), .partial_sum_in12(reg_psum14_5_2), .weight_in11(reg_weight14_5_1), .weight_in12(reg_weight14_5_2), .activation_in11(reg_activation15_4_1), .activation_in21(reg_activation15_4_2), .reg_partial_sum21(reg_psum15_5_1), .reg_partial_sum22(reg_psum15_5_2), .reg_weight21(reg_weight15_5_1), .reg_weight22(reg_weight15_5_2), .reg_activation12(reg_activation15_5_1), .reg_activation22(reg_activation15_5_2), .weight_en(weight_en));
SA22 U15_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_6_1), .partial_sum_in12(reg_psum14_6_2), .weight_in11(reg_weight14_6_1), .weight_in12(reg_weight14_6_2), .activation_in11(reg_activation15_5_1), .activation_in21(reg_activation15_5_2), .reg_partial_sum21(reg_psum15_6_1), .reg_partial_sum22(reg_psum15_6_2), .reg_weight21(reg_weight15_6_1), .reg_weight22(reg_weight15_6_2), .reg_activation12(reg_activation15_6_1), .reg_activation22(reg_activation15_6_2), .weight_en(weight_en));
SA22 U15_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_7_1), .partial_sum_in12(reg_psum14_7_2), .weight_in11(reg_weight14_7_1), .weight_in12(reg_weight14_7_2), .activation_in11(reg_activation15_6_1), .activation_in21(reg_activation15_6_2), .reg_partial_sum21(reg_psum15_7_1), .reg_partial_sum22(reg_psum15_7_2), .reg_weight21(reg_weight15_7_1), .reg_weight22(reg_weight15_7_2), .reg_activation12(reg_activation15_7_1), .reg_activation22(reg_activation15_7_2), .weight_en(weight_en));
SA22 U15_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_8_1), .partial_sum_in12(reg_psum14_8_2), .weight_in11(reg_weight14_8_1), .weight_in12(reg_weight14_8_2), .activation_in11(reg_activation15_7_1), .activation_in21(reg_activation15_7_2), .reg_partial_sum21(reg_psum15_8_1), .reg_partial_sum22(reg_psum15_8_2), .reg_weight21(reg_weight15_8_1), .reg_weight22(reg_weight15_8_2), .reg_activation12(reg_activation15_8_1), .reg_activation22(reg_activation15_8_2), .weight_en(weight_en));
SA22 U15_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_9_1), .partial_sum_in12(reg_psum14_9_2), .weight_in11(reg_weight14_9_1), .weight_in12(reg_weight14_9_2), .activation_in11(reg_activation15_8_1), .activation_in21(reg_activation15_8_2), .reg_partial_sum21(reg_psum15_9_1), .reg_partial_sum22(reg_psum15_9_2), .reg_weight21(reg_weight15_9_1), .reg_weight22(reg_weight15_9_2), .reg_activation12(reg_activation15_9_1), .reg_activation22(reg_activation15_9_2), .weight_en(weight_en));
SA22 U15_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_10_1), .partial_sum_in12(reg_psum14_10_2), .weight_in11(reg_weight14_10_1), .weight_in12(reg_weight14_10_2), .activation_in11(reg_activation15_9_1), .activation_in21(reg_activation15_9_2), .reg_partial_sum21(reg_psum15_10_1), .reg_partial_sum22(reg_psum15_10_2), .reg_weight21(reg_weight15_10_1), .reg_weight22(reg_weight15_10_2), .reg_activation12(reg_activation15_10_1), .reg_activation22(reg_activation15_10_2), .weight_en(weight_en));
SA22 U15_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_11_1), .partial_sum_in12(reg_psum14_11_2), .weight_in11(reg_weight14_11_1), .weight_in12(reg_weight14_11_2), .activation_in11(reg_activation15_10_1), .activation_in21(reg_activation15_10_2), .reg_partial_sum21(reg_psum15_11_1), .reg_partial_sum22(reg_psum15_11_2), .reg_weight21(reg_weight15_11_1), .reg_weight22(reg_weight15_11_2), .reg_activation12(reg_activation15_11_1), .reg_activation22(reg_activation15_11_2), .weight_en(weight_en));
SA22 U15_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_12_1), .partial_sum_in12(reg_psum14_12_2), .weight_in11(reg_weight14_12_1), .weight_in12(reg_weight14_12_2), .activation_in11(reg_activation15_11_1), .activation_in21(reg_activation15_11_2), .reg_partial_sum21(reg_psum15_12_1), .reg_partial_sum22(reg_psum15_12_2), .reg_weight21(reg_weight15_12_1), .reg_weight22(reg_weight15_12_2), .reg_activation12(reg_activation15_12_1), .reg_activation22(reg_activation15_12_2), .weight_en(weight_en));
SA22 U15_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_13_1), .partial_sum_in12(reg_psum14_13_2), .weight_in11(reg_weight14_13_1), .weight_in12(reg_weight14_13_2), .activation_in11(reg_activation15_12_1), .activation_in21(reg_activation15_12_2), .reg_partial_sum21(reg_psum15_13_1), .reg_partial_sum22(reg_psum15_13_2), .reg_weight21(reg_weight15_13_1), .reg_weight22(reg_weight15_13_2), .reg_activation12(reg_activation15_13_1), .reg_activation22(reg_activation15_13_2), .weight_en(weight_en));
SA22 U15_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_14_1), .partial_sum_in12(reg_psum14_14_2), .weight_in11(reg_weight14_14_1), .weight_in12(reg_weight14_14_2), .activation_in11(reg_activation15_13_1), .activation_in21(reg_activation15_13_2), .reg_partial_sum21(reg_psum15_14_1), .reg_partial_sum22(reg_psum15_14_2), .reg_weight21(reg_weight15_14_1), .reg_weight22(reg_weight15_14_2), .reg_activation12(reg_activation15_14_1), .reg_activation22(reg_activation15_14_2), .weight_en(weight_en));
SA22 U15_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_15_1), .partial_sum_in12(reg_psum14_15_2), .weight_in11(reg_weight14_15_1), .weight_in12(reg_weight14_15_2), .activation_in11(reg_activation15_14_1), .activation_in21(reg_activation15_14_2), .reg_partial_sum21(reg_psum15_15_1), .reg_partial_sum22(reg_psum15_15_2), .reg_weight21(reg_weight15_15_1), .reg_weight22(reg_weight15_15_2), .reg_activation12(reg_activation15_15_1), .reg_activation22(reg_activation15_15_2), .weight_en(weight_en));
SA22 U15_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_16_1), .partial_sum_in12(reg_psum14_16_2), .weight_in11(reg_weight14_16_1), .weight_in12(reg_weight14_16_2), .activation_in11(reg_activation15_15_1), .activation_in21(reg_activation15_15_2), .reg_partial_sum21(reg_psum15_16_1), .reg_partial_sum22(reg_psum15_16_2), .reg_weight21(reg_weight15_16_1), .reg_weight22(reg_weight15_16_2), .reg_activation12(reg_activation15_16_1), .reg_activation22(reg_activation15_16_2), .weight_en(weight_en));
SA22 U15_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_17_1), .partial_sum_in12(reg_psum14_17_2), .weight_in11(reg_weight14_17_1), .weight_in12(reg_weight14_17_2), .activation_in11(reg_activation15_16_1), .activation_in21(reg_activation15_16_2), .reg_partial_sum21(reg_psum15_17_1), .reg_partial_sum22(reg_psum15_17_2), .reg_weight21(reg_weight15_17_1), .reg_weight22(reg_weight15_17_2), .reg_activation12(reg_activation15_17_1), .reg_activation22(reg_activation15_17_2), .weight_en(weight_en));
SA22 U15_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_18_1), .partial_sum_in12(reg_psum14_18_2), .weight_in11(reg_weight14_18_1), .weight_in12(reg_weight14_18_2), .activation_in11(reg_activation15_17_1), .activation_in21(reg_activation15_17_2), .reg_partial_sum21(reg_psum15_18_1), .reg_partial_sum22(reg_psum15_18_2), .reg_weight21(reg_weight15_18_1), .reg_weight22(reg_weight15_18_2), .reg_activation12(reg_activation15_18_1), .reg_activation22(reg_activation15_18_2), .weight_en(weight_en));
SA22 U15_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_19_1), .partial_sum_in12(reg_psum14_19_2), .weight_in11(reg_weight14_19_1), .weight_in12(reg_weight14_19_2), .activation_in11(reg_activation15_18_1), .activation_in21(reg_activation15_18_2), .reg_partial_sum21(reg_psum15_19_1), .reg_partial_sum22(reg_psum15_19_2), .reg_weight21(reg_weight15_19_1), .reg_weight22(reg_weight15_19_2), .reg_activation12(reg_activation15_19_1), .reg_activation22(reg_activation15_19_2), .weight_en(weight_en));
SA22 U15_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_20_1), .partial_sum_in12(reg_psum14_20_2), .weight_in11(reg_weight14_20_1), .weight_in12(reg_weight14_20_2), .activation_in11(reg_activation15_19_1), .activation_in21(reg_activation15_19_2), .reg_partial_sum21(reg_psum15_20_1), .reg_partial_sum22(reg_psum15_20_2), .reg_weight21(reg_weight15_20_1), .reg_weight22(reg_weight15_20_2), .reg_activation12(reg_activation15_20_1), .reg_activation22(reg_activation15_20_2), .weight_en(weight_en));
SA22 U15_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_21_1), .partial_sum_in12(reg_psum14_21_2), .weight_in11(reg_weight14_21_1), .weight_in12(reg_weight14_21_2), .activation_in11(reg_activation15_20_1), .activation_in21(reg_activation15_20_2), .reg_partial_sum21(reg_psum15_21_1), .reg_partial_sum22(reg_psum15_21_2), .reg_weight21(reg_weight15_21_1), .reg_weight22(reg_weight15_21_2), .reg_activation12(reg_activation15_21_1), .reg_activation22(reg_activation15_21_2), .weight_en(weight_en));
SA22 U15_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_22_1), .partial_sum_in12(reg_psum14_22_2), .weight_in11(reg_weight14_22_1), .weight_in12(reg_weight14_22_2), .activation_in11(reg_activation15_21_1), .activation_in21(reg_activation15_21_2), .reg_partial_sum21(reg_psum15_22_1), .reg_partial_sum22(reg_psum15_22_2), .reg_weight21(reg_weight15_22_1), .reg_weight22(reg_weight15_22_2), .reg_activation12(reg_activation15_22_1), .reg_activation22(reg_activation15_22_2), .weight_en(weight_en));
SA22 U15_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_23_1), .partial_sum_in12(reg_psum14_23_2), .weight_in11(reg_weight14_23_1), .weight_in12(reg_weight14_23_2), .activation_in11(reg_activation15_22_1), .activation_in21(reg_activation15_22_2), .reg_partial_sum21(reg_psum15_23_1), .reg_partial_sum22(reg_psum15_23_2), .reg_weight21(reg_weight15_23_1), .reg_weight22(reg_weight15_23_2), .reg_activation12(reg_activation15_23_1), .reg_activation22(reg_activation15_23_2), .weight_en(weight_en));
SA22 U15_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_24_1), .partial_sum_in12(reg_psum14_24_2), .weight_in11(reg_weight14_24_1), .weight_in12(reg_weight14_24_2), .activation_in11(reg_activation15_23_1), .activation_in21(reg_activation15_23_2), .reg_partial_sum21(reg_psum15_24_1), .reg_partial_sum22(reg_psum15_24_2), .reg_weight21(reg_weight15_24_1), .reg_weight22(reg_weight15_24_2), .reg_activation12(reg_activation15_24_1), .reg_activation22(reg_activation15_24_2), .weight_en(weight_en));
SA22 U15_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_25_1), .partial_sum_in12(reg_psum14_25_2), .weight_in11(reg_weight14_25_1), .weight_in12(reg_weight14_25_2), .activation_in11(reg_activation15_24_1), .activation_in21(reg_activation15_24_2), .reg_partial_sum21(reg_psum15_25_1), .reg_partial_sum22(reg_psum15_25_2), .reg_weight21(reg_weight15_25_1), .reg_weight22(reg_weight15_25_2), .reg_activation12(reg_activation15_25_1), .reg_activation22(reg_activation15_25_2), .weight_en(weight_en));
SA22 U15_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_26_1), .partial_sum_in12(reg_psum14_26_2), .weight_in11(reg_weight14_26_1), .weight_in12(reg_weight14_26_2), .activation_in11(reg_activation15_25_1), .activation_in21(reg_activation15_25_2), .reg_partial_sum21(reg_psum15_26_1), .reg_partial_sum22(reg_psum15_26_2), .reg_weight21(reg_weight15_26_1), .reg_weight22(reg_weight15_26_2), .reg_activation12(reg_activation15_26_1), .reg_activation22(reg_activation15_26_2), .weight_en(weight_en));
SA22 U15_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_27_1), .partial_sum_in12(reg_psum14_27_2), .weight_in11(reg_weight14_27_1), .weight_in12(reg_weight14_27_2), .activation_in11(reg_activation15_26_1), .activation_in21(reg_activation15_26_2), .reg_partial_sum21(reg_psum15_27_1), .reg_partial_sum22(reg_psum15_27_2), .reg_weight21(reg_weight15_27_1), .reg_weight22(reg_weight15_27_2), .reg_activation12(reg_activation15_27_1), .reg_activation22(reg_activation15_27_2), .weight_en(weight_en));
SA22 U15_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_28_1), .partial_sum_in12(reg_psum14_28_2), .weight_in11(reg_weight14_28_1), .weight_in12(reg_weight14_28_2), .activation_in11(reg_activation15_27_1), .activation_in21(reg_activation15_27_2), .reg_partial_sum21(reg_psum15_28_1), .reg_partial_sum22(reg_psum15_28_2), .reg_weight21(reg_weight15_28_1), .reg_weight22(reg_weight15_28_2), .reg_activation12(reg_activation15_28_1), .reg_activation22(reg_activation15_28_2), .weight_en(weight_en));
SA22 U15_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_29_1), .partial_sum_in12(reg_psum14_29_2), .weight_in11(reg_weight14_29_1), .weight_in12(reg_weight14_29_2), .activation_in11(reg_activation15_28_1), .activation_in21(reg_activation15_28_2), .reg_partial_sum21(reg_psum15_29_1), .reg_partial_sum22(reg_psum15_29_2), .reg_weight21(reg_weight15_29_1), .reg_weight22(reg_weight15_29_2), .reg_activation12(reg_activation15_29_1), .reg_activation22(reg_activation15_29_2), .weight_en(weight_en));
SA22 U15_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_30_1), .partial_sum_in12(reg_psum14_30_2), .weight_in11(reg_weight14_30_1), .weight_in12(reg_weight14_30_2), .activation_in11(reg_activation15_29_1), .activation_in21(reg_activation15_29_2), .reg_partial_sum21(reg_psum15_30_1), .reg_partial_sum22(reg_psum15_30_2), .reg_weight21(reg_weight15_30_1), .reg_weight22(reg_weight15_30_2), .reg_activation12(reg_activation15_30_1), .reg_activation22(reg_activation15_30_2), .weight_en(weight_en));
SA22 U15_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_31_1), .partial_sum_in12(reg_psum14_31_2), .weight_in11(reg_weight14_31_1), .weight_in12(reg_weight14_31_2), .activation_in11(reg_activation15_30_1), .activation_in21(reg_activation15_30_2), .reg_partial_sum21(reg_psum15_31_1), .reg_partial_sum22(reg_psum15_31_2), .reg_weight21(reg_weight15_31_1), .reg_weight22(reg_weight15_31_2), .reg_activation12(reg_activation15_31_1), .reg_activation22(reg_activation15_31_2), .weight_en(weight_en));
SA22 U15_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum14_32_1), .partial_sum_in12(reg_psum14_32_2), .weight_in11(reg_weight14_32_1), .weight_in12(reg_weight14_32_2), .activation_in11(reg_activation15_31_1), .activation_in21(reg_activation15_31_2), .reg_partial_sum21(reg_psum15_32_1), .reg_partial_sum22(reg_psum15_32_2), .reg_weight21(reg_weight15_32_1), .reg_weight22(reg_weight15_32_2), .weight_en(weight_en));
SA22 U16_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_1_1), .partial_sum_in12(reg_psum15_1_2), .weight_in11(reg_weight15_1_1), .weight_in12(reg_weight15_1_2), .activation_in11(in_activation16_1_1), .activation_in21(in_activation16_1_2), .reg_partial_sum21(reg_psum16_1_1), .reg_partial_sum22(reg_psum16_1_2), .reg_weight21(reg_weight16_1_1), .reg_weight22(reg_weight16_1_2), .reg_activation12(reg_activation16_1_1), .reg_activation22(reg_activation16_1_2), .weight_en(weight_en));
SA22 U16_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_2_1), .partial_sum_in12(reg_psum15_2_2), .weight_in11(reg_weight15_2_1), .weight_in12(reg_weight15_2_2), .activation_in11(reg_activation16_1_1), .activation_in21(reg_activation16_1_2), .reg_partial_sum21(reg_psum16_2_1), .reg_partial_sum22(reg_psum16_2_2), .reg_weight21(reg_weight16_2_1), .reg_weight22(reg_weight16_2_2), .reg_activation12(reg_activation16_2_1), .reg_activation22(reg_activation16_2_2), .weight_en(weight_en));
SA22 U16_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_3_1), .partial_sum_in12(reg_psum15_3_2), .weight_in11(reg_weight15_3_1), .weight_in12(reg_weight15_3_2), .activation_in11(reg_activation16_2_1), .activation_in21(reg_activation16_2_2), .reg_partial_sum21(reg_psum16_3_1), .reg_partial_sum22(reg_psum16_3_2), .reg_weight21(reg_weight16_3_1), .reg_weight22(reg_weight16_3_2), .reg_activation12(reg_activation16_3_1), .reg_activation22(reg_activation16_3_2), .weight_en(weight_en));
SA22 U16_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_4_1), .partial_sum_in12(reg_psum15_4_2), .weight_in11(reg_weight15_4_1), .weight_in12(reg_weight15_4_2), .activation_in11(reg_activation16_3_1), .activation_in21(reg_activation16_3_2), .reg_partial_sum21(reg_psum16_4_1), .reg_partial_sum22(reg_psum16_4_2), .reg_weight21(reg_weight16_4_1), .reg_weight22(reg_weight16_4_2), .reg_activation12(reg_activation16_4_1), .reg_activation22(reg_activation16_4_2), .weight_en(weight_en));
SA22 U16_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_5_1), .partial_sum_in12(reg_psum15_5_2), .weight_in11(reg_weight15_5_1), .weight_in12(reg_weight15_5_2), .activation_in11(reg_activation16_4_1), .activation_in21(reg_activation16_4_2), .reg_partial_sum21(reg_psum16_5_1), .reg_partial_sum22(reg_psum16_5_2), .reg_weight21(reg_weight16_5_1), .reg_weight22(reg_weight16_5_2), .reg_activation12(reg_activation16_5_1), .reg_activation22(reg_activation16_5_2), .weight_en(weight_en));
SA22 U16_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_6_1), .partial_sum_in12(reg_psum15_6_2), .weight_in11(reg_weight15_6_1), .weight_in12(reg_weight15_6_2), .activation_in11(reg_activation16_5_1), .activation_in21(reg_activation16_5_2), .reg_partial_sum21(reg_psum16_6_1), .reg_partial_sum22(reg_psum16_6_2), .reg_weight21(reg_weight16_6_1), .reg_weight22(reg_weight16_6_2), .reg_activation12(reg_activation16_6_1), .reg_activation22(reg_activation16_6_2), .weight_en(weight_en));
SA22 U16_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_7_1), .partial_sum_in12(reg_psum15_7_2), .weight_in11(reg_weight15_7_1), .weight_in12(reg_weight15_7_2), .activation_in11(reg_activation16_6_1), .activation_in21(reg_activation16_6_2), .reg_partial_sum21(reg_psum16_7_1), .reg_partial_sum22(reg_psum16_7_2), .reg_weight21(reg_weight16_7_1), .reg_weight22(reg_weight16_7_2), .reg_activation12(reg_activation16_7_1), .reg_activation22(reg_activation16_7_2), .weight_en(weight_en));
SA22 U16_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_8_1), .partial_sum_in12(reg_psum15_8_2), .weight_in11(reg_weight15_8_1), .weight_in12(reg_weight15_8_2), .activation_in11(reg_activation16_7_1), .activation_in21(reg_activation16_7_2), .reg_partial_sum21(reg_psum16_8_1), .reg_partial_sum22(reg_psum16_8_2), .reg_weight21(reg_weight16_8_1), .reg_weight22(reg_weight16_8_2), .reg_activation12(reg_activation16_8_1), .reg_activation22(reg_activation16_8_2), .weight_en(weight_en));
SA22 U16_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_9_1), .partial_sum_in12(reg_psum15_9_2), .weight_in11(reg_weight15_9_1), .weight_in12(reg_weight15_9_2), .activation_in11(reg_activation16_8_1), .activation_in21(reg_activation16_8_2), .reg_partial_sum21(reg_psum16_9_1), .reg_partial_sum22(reg_psum16_9_2), .reg_weight21(reg_weight16_9_1), .reg_weight22(reg_weight16_9_2), .reg_activation12(reg_activation16_9_1), .reg_activation22(reg_activation16_9_2), .weight_en(weight_en));
SA22 U16_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_10_1), .partial_sum_in12(reg_psum15_10_2), .weight_in11(reg_weight15_10_1), .weight_in12(reg_weight15_10_2), .activation_in11(reg_activation16_9_1), .activation_in21(reg_activation16_9_2), .reg_partial_sum21(reg_psum16_10_1), .reg_partial_sum22(reg_psum16_10_2), .reg_weight21(reg_weight16_10_1), .reg_weight22(reg_weight16_10_2), .reg_activation12(reg_activation16_10_1), .reg_activation22(reg_activation16_10_2), .weight_en(weight_en));
SA22 U16_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_11_1), .partial_sum_in12(reg_psum15_11_2), .weight_in11(reg_weight15_11_1), .weight_in12(reg_weight15_11_2), .activation_in11(reg_activation16_10_1), .activation_in21(reg_activation16_10_2), .reg_partial_sum21(reg_psum16_11_1), .reg_partial_sum22(reg_psum16_11_2), .reg_weight21(reg_weight16_11_1), .reg_weight22(reg_weight16_11_2), .reg_activation12(reg_activation16_11_1), .reg_activation22(reg_activation16_11_2), .weight_en(weight_en));
SA22 U16_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_12_1), .partial_sum_in12(reg_psum15_12_2), .weight_in11(reg_weight15_12_1), .weight_in12(reg_weight15_12_2), .activation_in11(reg_activation16_11_1), .activation_in21(reg_activation16_11_2), .reg_partial_sum21(reg_psum16_12_1), .reg_partial_sum22(reg_psum16_12_2), .reg_weight21(reg_weight16_12_1), .reg_weight22(reg_weight16_12_2), .reg_activation12(reg_activation16_12_1), .reg_activation22(reg_activation16_12_2), .weight_en(weight_en));
SA22 U16_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_13_1), .partial_sum_in12(reg_psum15_13_2), .weight_in11(reg_weight15_13_1), .weight_in12(reg_weight15_13_2), .activation_in11(reg_activation16_12_1), .activation_in21(reg_activation16_12_2), .reg_partial_sum21(reg_psum16_13_1), .reg_partial_sum22(reg_psum16_13_2), .reg_weight21(reg_weight16_13_1), .reg_weight22(reg_weight16_13_2), .reg_activation12(reg_activation16_13_1), .reg_activation22(reg_activation16_13_2), .weight_en(weight_en));
SA22 U16_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_14_1), .partial_sum_in12(reg_psum15_14_2), .weight_in11(reg_weight15_14_1), .weight_in12(reg_weight15_14_2), .activation_in11(reg_activation16_13_1), .activation_in21(reg_activation16_13_2), .reg_partial_sum21(reg_psum16_14_1), .reg_partial_sum22(reg_psum16_14_2), .reg_weight21(reg_weight16_14_1), .reg_weight22(reg_weight16_14_2), .reg_activation12(reg_activation16_14_1), .reg_activation22(reg_activation16_14_2), .weight_en(weight_en));
SA22 U16_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_15_1), .partial_sum_in12(reg_psum15_15_2), .weight_in11(reg_weight15_15_1), .weight_in12(reg_weight15_15_2), .activation_in11(reg_activation16_14_1), .activation_in21(reg_activation16_14_2), .reg_partial_sum21(reg_psum16_15_1), .reg_partial_sum22(reg_psum16_15_2), .reg_weight21(reg_weight16_15_1), .reg_weight22(reg_weight16_15_2), .reg_activation12(reg_activation16_15_1), .reg_activation22(reg_activation16_15_2), .weight_en(weight_en));
SA22 U16_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_16_1), .partial_sum_in12(reg_psum15_16_2), .weight_in11(reg_weight15_16_1), .weight_in12(reg_weight15_16_2), .activation_in11(reg_activation16_15_1), .activation_in21(reg_activation16_15_2), .reg_partial_sum21(reg_psum16_16_1), .reg_partial_sum22(reg_psum16_16_2), .reg_weight21(reg_weight16_16_1), .reg_weight22(reg_weight16_16_2), .reg_activation12(reg_activation16_16_1), .reg_activation22(reg_activation16_16_2), .weight_en(weight_en));
SA22 U16_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_17_1), .partial_sum_in12(reg_psum15_17_2), .weight_in11(reg_weight15_17_1), .weight_in12(reg_weight15_17_2), .activation_in11(reg_activation16_16_1), .activation_in21(reg_activation16_16_2), .reg_partial_sum21(reg_psum16_17_1), .reg_partial_sum22(reg_psum16_17_2), .reg_weight21(reg_weight16_17_1), .reg_weight22(reg_weight16_17_2), .reg_activation12(reg_activation16_17_1), .reg_activation22(reg_activation16_17_2), .weight_en(weight_en));
SA22 U16_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_18_1), .partial_sum_in12(reg_psum15_18_2), .weight_in11(reg_weight15_18_1), .weight_in12(reg_weight15_18_2), .activation_in11(reg_activation16_17_1), .activation_in21(reg_activation16_17_2), .reg_partial_sum21(reg_psum16_18_1), .reg_partial_sum22(reg_psum16_18_2), .reg_weight21(reg_weight16_18_1), .reg_weight22(reg_weight16_18_2), .reg_activation12(reg_activation16_18_1), .reg_activation22(reg_activation16_18_2), .weight_en(weight_en));
SA22 U16_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_19_1), .partial_sum_in12(reg_psum15_19_2), .weight_in11(reg_weight15_19_1), .weight_in12(reg_weight15_19_2), .activation_in11(reg_activation16_18_1), .activation_in21(reg_activation16_18_2), .reg_partial_sum21(reg_psum16_19_1), .reg_partial_sum22(reg_psum16_19_2), .reg_weight21(reg_weight16_19_1), .reg_weight22(reg_weight16_19_2), .reg_activation12(reg_activation16_19_1), .reg_activation22(reg_activation16_19_2), .weight_en(weight_en));
SA22 U16_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_20_1), .partial_sum_in12(reg_psum15_20_2), .weight_in11(reg_weight15_20_1), .weight_in12(reg_weight15_20_2), .activation_in11(reg_activation16_19_1), .activation_in21(reg_activation16_19_2), .reg_partial_sum21(reg_psum16_20_1), .reg_partial_sum22(reg_psum16_20_2), .reg_weight21(reg_weight16_20_1), .reg_weight22(reg_weight16_20_2), .reg_activation12(reg_activation16_20_1), .reg_activation22(reg_activation16_20_2), .weight_en(weight_en));
SA22 U16_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_21_1), .partial_sum_in12(reg_psum15_21_2), .weight_in11(reg_weight15_21_1), .weight_in12(reg_weight15_21_2), .activation_in11(reg_activation16_20_1), .activation_in21(reg_activation16_20_2), .reg_partial_sum21(reg_psum16_21_1), .reg_partial_sum22(reg_psum16_21_2), .reg_weight21(reg_weight16_21_1), .reg_weight22(reg_weight16_21_2), .reg_activation12(reg_activation16_21_1), .reg_activation22(reg_activation16_21_2), .weight_en(weight_en));
SA22 U16_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_22_1), .partial_sum_in12(reg_psum15_22_2), .weight_in11(reg_weight15_22_1), .weight_in12(reg_weight15_22_2), .activation_in11(reg_activation16_21_1), .activation_in21(reg_activation16_21_2), .reg_partial_sum21(reg_psum16_22_1), .reg_partial_sum22(reg_psum16_22_2), .reg_weight21(reg_weight16_22_1), .reg_weight22(reg_weight16_22_2), .reg_activation12(reg_activation16_22_1), .reg_activation22(reg_activation16_22_2), .weight_en(weight_en));
SA22 U16_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_23_1), .partial_sum_in12(reg_psum15_23_2), .weight_in11(reg_weight15_23_1), .weight_in12(reg_weight15_23_2), .activation_in11(reg_activation16_22_1), .activation_in21(reg_activation16_22_2), .reg_partial_sum21(reg_psum16_23_1), .reg_partial_sum22(reg_psum16_23_2), .reg_weight21(reg_weight16_23_1), .reg_weight22(reg_weight16_23_2), .reg_activation12(reg_activation16_23_1), .reg_activation22(reg_activation16_23_2), .weight_en(weight_en));
SA22 U16_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_24_1), .partial_sum_in12(reg_psum15_24_2), .weight_in11(reg_weight15_24_1), .weight_in12(reg_weight15_24_2), .activation_in11(reg_activation16_23_1), .activation_in21(reg_activation16_23_2), .reg_partial_sum21(reg_psum16_24_1), .reg_partial_sum22(reg_psum16_24_2), .reg_weight21(reg_weight16_24_1), .reg_weight22(reg_weight16_24_2), .reg_activation12(reg_activation16_24_1), .reg_activation22(reg_activation16_24_2), .weight_en(weight_en));
SA22 U16_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_25_1), .partial_sum_in12(reg_psum15_25_2), .weight_in11(reg_weight15_25_1), .weight_in12(reg_weight15_25_2), .activation_in11(reg_activation16_24_1), .activation_in21(reg_activation16_24_2), .reg_partial_sum21(reg_psum16_25_1), .reg_partial_sum22(reg_psum16_25_2), .reg_weight21(reg_weight16_25_1), .reg_weight22(reg_weight16_25_2), .reg_activation12(reg_activation16_25_1), .reg_activation22(reg_activation16_25_2), .weight_en(weight_en));
SA22 U16_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_26_1), .partial_sum_in12(reg_psum15_26_2), .weight_in11(reg_weight15_26_1), .weight_in12(reg_weight15_26_2), .activation_in11(reg_activation16_25_1), .activation_in21(reg_activation16_25_2), .reg_partial_sum21(reg_psum16_26_1), .reg_partial_sum22(reg_psum16_26_2), .reg_weight21(reg_weight16_26_1), .reg_weight22(reg_weight16_26_2), .reg_activation12(reg_activation16_26_1), .reg_activation22(reg_activation16_26_2), .weight_en(weight_en));
SA22 U16_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_27_1), .partial_sum_in12(reg_psum15_27_2), .weight_in11(reg_weight15_27_1), .weight_in12(reg_weight15_27_2), .activation_in11(reg_activation16_26_1), .activation_in21(reg_activation16_26_2), .reg_partial_sum21(reg_psum16_27_1), .reg_partial_sum22(reg_psum16_27_2), .reg_weight21(reg_weight16_27_1), .reg_weight22(reg_weight16_27_2), .reg_activation12(reg_activation16_27_1), .reg_activation22(reg_activation16_27_2), .weight_en(weight_en));
SA22 U16_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_28_1), .partial_sum_in12(reg_psum15_28_2), .weight_in11(reg_weight15_28_1), .weight_in12(reg_weight15_28_2), .activation_in11(reg_activation16_27_1), .activation_in21(reg_activation16_27_2), .reg_partial_sum21(reg_psum16_28_1), .reg_partial_sum22(reg_psum16_28_2), .reg_weight21(reg_weight16_28_1), .reg_weight22(reg_weight16_28_2), .reg_activation12(reg_activation16_28_1), .reg_activation22(reg_activation16_28_2), .weight_en(weight_en));
SA22 U16_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_29_1), .partial_sum_in12(reg_psum15_29_2), .weight_in11(reg_weight15_29_1), .weight_in12(reg_weight15_29_2), .activation_in11(reg_activation16_28_1), .activation_in21(reg_activation16_28_2), .reg_partial_sum21(reg_psum16_29_1), .reg_partial_sum22(reg_psum16_29_2), .reg_weight21(reg_weight16_29_1), .reg_weight22(reg_weight16_29_2), .reg_activation12(reg_activation16_29_1), .reg_activation22(reg_activation16_29_2), .weight_en(weight_en));
SA22 U16_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_30_1), .partial_sum_in12(reg_psum15_30_2), .weight_in11(reg_weight15_30_1), .weight_in12(reg_weight15_30_2), .activation_in11(reg_activation16_29_1), .activation_in21(reg_activation16_29_2), .reg_partial_sum21(reg_psum16_30_1), .reg_partial_sum22(reg_psum16_30_2), .reg_weight21(reg_weight16_30_1), .reg_weight22(reg_weight16_30_2), .reg_activation12(reg_activation16_30_1), .reg_activation22(reg_activation16_30_2), .weight_en(weight_en));
SA22 U16_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_31_1), .partial_sum_in12(reg_psum15_31_2), .weight_in11(reg_weight15_31_1), .weight_in12(reg_weight15_31_2), .activation_in11(reg_activation16_30_1), .activation_in21(reg_activation16_30_2), .reg_partial_sum21(reg_psum16_31_1), .reg_partial_sum22(reg_psum16_31_2), .reg_weight21(reg_weight16_31_1), .reg_weight22(reg_weight16_31_2), .reg_activation12(reg_activation16_31_1), .reg_activation22(reg_activation16_31_2), .weight_en(weight_en));
SA22 U16_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum15_32_1), .partial_sum_in12(reg_psum15_32_2), .weight_in11(reg_weight15_32_1), .weight_in12(reg_weight15_32_2), .activation_in11(reg_activation16_31_1), .activation_in21(reg_activation16_31_2), .reg_partial_sum21(reg_psum16_32_1), .reg_partial_sum22(reg_psum16_32_2), .reg_weight21(reg_weight16_32_1), .reg_weight22(reg_weight16_32_2), .weight_en(weight_en));
SA22 U17_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_1_1), .partial_sum_in12(reg_psum16_1_2), .weight_in11(reg_weight16_1_1), .weight_in12(reg_weight16_1_2), .activation_in11(in_activation17_1_1), .activation_in21(in_activation17_1_2), .reg_partial_sum21(reg_psum17_1_1), .reg_partial_sum22(reg_psum17_1_2), .reg_weight21(reg_weight17_1_1), .reg_weight22(reg_weight17_1_2), .reg_activation12(reg_activation17_1_1), .reg_activation22(reg_activation17_1_2), .weight_en(weight_en));
SA22 U17_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_2_1), .partial_sum_in12(reg_psum16_2_2), .weight_in11(reg_weight16_2_1), .weight_in12(reg_weight16_2_2), .activation_in11(reg_activation17_1_1), .activation_in21(reg_activation17_1_2), .reg_partial_sum21(reg_psum17_2_1), .reg_partial_sum22(reg_psum17_2_2), .reg_weight21(reg_weight17_2_1), .reg_weight22(reg_weight17_2_2), .reg_activation12(reg_activation17_2_1), .reg_activation22(reg_activation17_2_2), .weight_en(weight_en));
SA22 U17_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_3_1), .partial_sum_in12(reg_psum16_3_2), .weight_in11(reg_weight16_3_1), .weight_in12(reg_weight16_3_2), .activation_in11(reg_activation17_2_1), .activation_in21(reg_activation17_2_2), .reg_partial_sum21(reg_psum17_3_1), .reg_partial_sum22(reg_psum17_3_2), .reg_weight21(reg_weight17_3_1), .reg_weight22(reg_weight17_3_2), .reg_activation12(reg_activation17_3_1), .reg_activation22(reg_activation17_3_2), .weight_en(weight_en));
SA22 U17_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_4_1), .partial_sum_in12(reg_psum16_4_2), .weight_in11(reg_weight16_4_1), .weight_in12(reg_weight16_4_2), .activation_in11(reg_activation17_3_1), .activation_in21(reg_activation17_3_2), .reg_partial_sum21(reg_psum17_4_1), .reg_partial_sum22(reg_psum17_4_2), .reg_weight21(reg_weight17_4_1), .reg_weight22(reg_weight17_4_2), .reg_activation12(reg_activation17_4_1), .reg_activation22(reg_activation17_4_2), .weight_en(weight_en));
SA22 U17_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_5_1), .partial_sum_in12(reg_psum16_5_2), .weight_in11(reg_weight16_5_1), .weight_in12(reg_weight16_5_2), .activation_in11(reg_activation17_4_1), .activation_in21(reg_activation17_4_2), .reg_partial_sum21(reg_psum17_5_1), .reg_partial_sum22(reg_psum17_5_2), .reg_weight21(reg_weight17_5_1), .reg_weight22(reg_weight17_5_2), .reg_activation12(reg_activation17_5_1), .reg_activation22(reg_activation17_5_2), .weight_en(weight_en));
SA22 U17_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_6_1), .partial_sum_in12(reg_psum16_6_2), .weight_in11(reg_weight16_6_1), .weight_in12(reg_weight16_6_2), .activation_in11(reg_activation17_5_1), .activation_in21(reg_activation17_5_2), .reg_partial_sum21(reg_psum17_6_1), .reg_partial_sum22(reg_psum17_6_2), .reg_weight21(reg_weight17_6_1), .reg_weight22(reg_weight17_6_2), .reg_activation12(reg_activation17_6_1), .reg_activation22(reg_activation17_6_2), .weight_en(weight_en));
SA22 U17_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_7_1), .partial_sum_in12(reg_psum16_7_2), .weight_in11(reg_weight16_7_1), .weight_in12(reg_weight16_7_2), .activation_in11(reg_activation17_6_1), .activation_in21(reg_activation17_6_2), .reg_partial_sum21(reg_psum17_7_1), .reg_partial_sum22(reg_psum17_7_2), .reg_weight21(reg_weight17_7_1), .reg_weight22(reg_weight17_7_2), .reg_activation12(reg_activation17_7_1), .reg_activation22(reg_activation17_7_2), .weight_en(weight_en));
SA22 U17_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_8_1), .partial_sum_in12(reg_psum16_8_2), .weight_in11(reg_weight16_8_1), .weight_in12(reg_weight16_8_2), .activation_in11(reg_activation17_7_1), .activation_in21(reg_activation17_7_2), .reg_partial_sum21(reg_psum17_8_1), .reg_partial_sum22(reg_psum17_8_2), .reg_weight21(reg_weight17_8_1), .reg_weight22(reg_weight17_8_2), .reg_activation12(reg_activation17_8_1), .reg_activation22(reg_activation17_8_2), .weight_en(weight_en));
SA22 U17_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_9_1), .partial_sum_in12(reg_psum16_9_2), .weight_in11(reg_weight16_9_1), .weight_in12(reg_weight16_9_2), .activation_in11(reg_activation17_8_1), .activation_in21(reg_activation17_8_2), .reg_partial_sum21(reg_psum17_9_1), .reg_partial_sum22(reg_psum17_9_2), .reg_weight21(reg_weight17_9_1), .reg_weight22(reg_weight17_9_2), .reg_activation12(reg_activation17_9_1), .reg_activation22(reg_activation17_9_2), .weight_en(weight_en));
SA22 U17_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_10_1), .partial_sum_in12(reg_psum16_10_2), .weight_in11(reg_weight16_10_1), .weight_in12(reg_weight16_10_2), .activation_in11(reg_activation17_9_1), .activation_in21(reg_activation17_9_2), .reg_partial_sum21(reg_psum17_10_1), .reg_partial_sum22(reg_psum17_10_2), .reg_weight21(reg_weight17_10_1), .reg_weight22(reg_weight17_10_2), .reg_activation12(reg_activation17_10_1), .reg_activation22(reg_activation17_10_2), .weight_en(weight_en));
SA22 U17_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_11_1), .partial_sum_in12(reg_psum16_11_2), .weight_in11(reg_weight16_11_1), .weight_in12(reg_weight16_11_2), .activation_in11(reg_activation17_10_1), .activation_in21(reg_activation17_10_2), .reg_partial_sum21(reg_psum17_11_1), .reg_partial_sum22(reg_psum17_11_2), .reg_weight21(reg_weight17_11_1), .reg_weight22(reg_weight17_11_2), .reg_activation12(reg_activation17_11_1), .reg_activation22(reg_activation17_11_2), .weight_en(weight_en));
SA22 U17_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_12_1), .partial_sum_in12(reg_psum16_12_2), .weight_in11(reg_weight16_12_1), .weight_in12(reg_weight16_12_2), .activation_in11(reg_activation17_11_1), .activation_in21(reg_activation17_11_2), .reg_partial_sum21(reg_psum17_12_1), .reg_partial_sum22(reg_psum17_12_2), .reg_weight21(reg_weight17_12_1), .reg_weight22(reg_weight17_12_2), .reg_activation12(reg_activation17_12_1), .reg_activation22(reg_activation17_12_2), .weight_en(weight_en));
SA22 U17_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_13_1), .partial_sum_in12(reg_psum16_13_2), .weight_in11(reg_weight16_13_1), .weight_in12(reg_weight16_13_2), .activation_in11(reg_activation17_12_1), .activation_in21(reg_activation17_12_2), .reg_partial_sum21(reg_psum17_13_1), .reg_partial_sum22(reg_psum17_13_2), .reg_weight21(reg_weight17_13_1), .reg_weight22(reg_weight17_13_2), .reg_activation12(reg_activation17_13_1), .reg_activation22(reg_activation17_13_2), .weight_en(weight_en));
SA22 U17_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_14_1), .partial_sum_in12(reg_psum16_14_2), .weight_in11(reg_weight16_14_1), .weight_in12(reg_weight16_14_2), .activation_in11(reg_activation17_13_1), .activation_in21(reg_activation17_13_2), .reg_partial_sum21(reg_psum17_14_1), .reg_partial_sum22(reg_psum17_14_2), .reg_weight21(reg_weight17_14_1), .reg_weight22(reg_weight17_14_2), .reg_activation12(reg_activation17_14_1), .reg_activation22(reg_activation17_14_2), .weight_en(weight_en));
SA22 U17_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_15_1), .partial_sum_in12(reg_psum16_15_2), .weight_in11(reg_weight16_15_1), .weight_in12(reg_weight16_15_2), .activation_in11(reg_activation17_14_1), .activation_in21(reg_activation17_14_2), .reg_partial_sum21(reg_psum17_15_1), .reg_partial_sum22(reg_psum17_15_2), .reg_weight21(reg_weight17_15_1), .reg_weight22(reg_weight17_15_2), .reg_activation12(reg_activation17_15_1), .reg_activation22(reg_activation17_15_2), .weight_en(weight_en));
SA22 U17_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_16_1), .partial_sum_in12(reg_psum16_16_2), .weight_in11(reg_weight16_16_1), .weight_in12(reg_weight16_16_2), .activation_in11(reg_activation17_15_1), .activation_in21(reg_activation17_15_2), .reg_partial_sum21(reg_psum17_16_1), .reg_partial_sum22(reg_psum17_16_2), .reg_weight21(reg_weight17_16_1), .reg_weight22(reg_weight17_16_2), .reg_activation12(reg_activation17_16_1), .reg_activation22(reg_activation17_16_2), .weight_en(weight_en));
SA22 U17_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_17_1), .partial_sum_in12(reg_psum16_17_2), .weight_in11(reg_weight16_17_1), .weight_in12(reg_weight16_17_2), .activation_in11(reg_activation17_16_1), .activation_in21(reg_activation17_16_2), .reg_partial_sum21(reg_psum17_17_1), .reg_partial_sum22(reg_psum17_17_2), .reg_weight21(reg_weight17_17_1), .reg_weight22(reg_weight17_17_2), .reg_activation12(reg_activation17_17_1), .reg_activation22(reg_activation17_17_2), .weight_en(weight_en));
SA22 U17_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_18_1), .partial_sum_in12(reg_psum16_18_2), .weight_in11(reg_weight16_18_1), .weight_in12(reg_weight16_18_2), .activation_in11(reg_activation17_17_1), .activation_in21(reg_activation17_17_2), .reg_partial_sum21(reg_psum17_18_1), .reg_partial_sum22(reg_psum17_18_2), .reg_weight21(reg_weight17_18_1), .reg_weight22(reg_weight17_18_2), .reg_activation12(reg_activation17_18_1), .reg_activation22(reg_activation17_18_2), .weight_en(weight_en));
SA22 U17_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_19_1), .partial_sum_in12(reg_psum16_19_2), .weight_in11(reg_weight16_19_1), .weight_in12(reg_weight16_19_2), .activation_in11(reg_activation17_18_1), .activation_in21(reg_activation17_18_2), .reg_partial_sum21(reg_psum17_19_1), .reg_partial_sum22(reg_psum17_19_2), .reg_weight21(reg_weight17_19_1), .reg_weight22(reg_weight17_19_2), .reg_activation12(reg_activation17_19_1), .reg_activation22(reg_activation17_19_2), .weight_en(weight_en));
SA22 U17_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_20_1), .partial_sum_in12(reg_psum16_20_2), .weight_in11(reg_weight16_20_1), .weight_in12(reg_weight16_20_2), .activation_in11(reg_activation17_19_1), .activation_in21(reg_activation17_19_2), .reg_partial_sum21(reg_psum17_20_1), .reg_partial_sum22(reg_psum17_20_2), .reg_weight21(reg_weight17_20_1), .reg_weight22(reg_weight17_20_2), .reg_activation12(reg_activation17_20_1), .reg_activation22(reg_activation17_20_2), .weight_en(weight_en));
SA22 U17_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_21_1), .partial_sum_in12(reg_psum16_21_2), .weight_in11(reg_weight16_21_1), .weight_in12(reg_weight16_21_2), .activation_in11(reg_activation17_20_1), .activation_in21(reg_activation17_20_2), .reg_partial_sum21(reg_psum17_21_1), .reg_partial_sum22(reg_psum17_21_2), .reg_weight21(reg_weight17_21_1), .reg_weight22(reg_weight17_21_2), .reg_activation12(reg_activation17_21_1), .reg_activation22(reg_activation17_21_2), .weight_en(weight_en));
SA22 U17_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_22_1), .partial_sum_in12(reg_psum16_22_2), .weight_in11(reg_weight16_22_1), .weight_in12(reg_weight16_22_2), .activation_in11(reg_activation17_21_1), .activation_in21(reg_activation17_21_2), .reg_partial_sum21(reg_psum17_22_1), .reg_partial_sum22(reg_psum17_22_2), .reg_weight21(reg_weight17_22_1), .reg_weight22(reg_weight17_22_2), .reg_activation12(reg_activation17_22_1), .reg_activation22(reg_activation17_22_2), .weight_en(weight_en));
SA22 U17_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_23_1), .partial_sum_in12(reg_psum16_23_2), .weight_in11(reg_weight16_23_1), .weight_in12(reg_weight16_23_2), .activation_in11(reg_activation17_22_1), .activation_in21(reg_activation17_22_2), .reg_partial_sum21(reg_psum17_23_1), .reg_partial_sum22(reg_psum17_23_2), .reg_weight21(reg_weight17_23_1), .reg_weight22(reg_weight17_23_2), .reg_activation12(reg_activation17_23_1), .reg_activation22(reg_activation17_23_2), .weight_en(weight_en));
SA22 U17_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_24_1), .partial_sum_in12(reg_psum16_24_2), .weight_in11(reg_weight16_24_1), .weight_in12(reg_weight16_24_2), .activation_in11(reg_activation17_23_1), .activation_in21(reg_activation17_23_2), .reg_partial_sum21(reg_psum17_24_1), .reg_partial_sum22(reg_psum17_24_2), .reg_weight21(reg_weight17_24_1), .reg_weight22(reg_weight17_24_2), .reg_activation12(reg_activation17_24_1), .reg_activation22(reg_activation17_24_2), .weight_en(weight_en));
SA22 U17_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_25_1), .partial_sum_in12(reg_psum16_25_2), .weight_in11(reg_weight16_25_1), .weight_in12(reg_weight16_25_2), .activation_in11(reg_activation17_24_1), .activation_in21(reg_activation17_24_2), .reg_partial_sum21(reg_psum17_25_1), .reg_partial_sum22(reg_psum17_25_2), .reg_weight21(reg_weight17_25_1), .reg_weight22(reg_weight17_25_2), .reg_activation12(reg_activation17_25_1), .reg_activation22(reg_activation17_25_2), .weight_en(weight_en));
SA22 U17_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_26_1), .partial_sum_in12(reg_psum16_26_2), .weight_in11(reg_weight16_26_1), .weight_in12(reg_weight16_26_2), .activation_in11(reg_activation17_25_1), .activation_in21(reg_activation17_25_2), .reg_partial_sum21(reg_psum17_26_1), .reg_partial_sum22(reg_psum17_26_2), .reg_weight21(reg_weight17_26_1), .reg_weight22(reg_weight17_26_2), .reg_activation12(reg_activation17_26_1), .reg_activation22(reg_activation17_26_2), .weight_en(weight_en));
SA22 U17_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_27_1), .partial_sum_in12(reg_psum16_27_2), .weight_in11(reg_weight16_27_1), .weight_in12(reg_weight16_27_2), .activation_in11(reg_activation17_26_1), .activation_in21(reg_activation17_26_2), .reg_partial_sum21(reg_psum17_27_1), .reg_partial_sum22(reg_psum17_27_2), .reg_weight21(reg_weight17_27_1), .reg_weight22(reg_weight17_27_2), .reg_activation12(reg_activation17_27_1), .reg_activation22(reg_activation17_27_2), .weight_en(weight_en));
SA22 U17_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_28_1), .partial_sum_in12(reg_psum16_28_2), .weight_in11(reg_weight16_28_1), .weight_in12(reg_weight16_28_2), .activation_in11(reg_activation17_27_1), .activation_in21(reg_activation17_27_2), .reg_partial_sum21(reg_psum17_28_1), .reg_partial_sum22(reg_psum17_28_2), .reg_weight21(reg_weight17_28_1), .reg_weight22(reg_weight17_28_2), .reg_activation12(reg_activation17_28_1), .reg_activation22(reg_activation17_28_2), .weight_en(weight_en));
SA22 U17_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_29_1), .partial_sum_in12(reg_psum16_29_2), .weight_in11(reg_weight16_29_1), .weight_in12(reg_weight16_29_2), .activation_in11(reg_activation17_28_1), .activation_in21(reg_activation17_28_2), .reg_partial_sum21(reg_psum17_29_1), .reg_partial_sum22(reg_psum17_29_2), .reg_weight21(reg_weight17_29_1), .reg_weight22(reg_weight17_29_2), .reg_activation12(reg_activation17_29_1), .reg_activation22(reg_activation17_29_2), .weight_en(weight_en));
SA22 U17_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_30_1), .partial_sum_in12(reg_psum16_30_2), .weight_in11(reg_weight16_30_1), .weight_in12(reg_weight16_30_2), .activation_in11(reg_activation17_29_1), .activation_in21(reg_activation17_29_2), .reg_partial_sum21(reg_psum17_30_1), .reg_partial_sum22(reg_psum17_30_2), .reg_weight21(reg_weight17_30_1), .reg_weight22(reg_weight17_30_2), .reg_activation12(reg_activation17_30_1), .reg_activation22(reg_activation17_30_2), .weight_en(weight_en));
SA22 U17_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_31_1), .partial_sum_in12(reg_psum16_31_2), .weight_in11(reg_weight16_31_1), .weight_in12(reg_weight16_31_2), .activation_in11(reg_activation17_30_1), .activation_in21(reg_activation17_30_2), .reg_partial_sum21(reg_psum17_31_1), .reg_partial_sum22(reg_psum17_31_2), .reg_weight21(reg_weight17_31_1), .reg_weight22(reg_weight17_31_2), .reg_activation12(reg_activation17_31_1), .reg_activation22(reg_activation17_31_2), .weight_en(weight_en));
SA22 U17_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum16_32_1), .partial_sum_in12(reg_psum16_32_2), .weight_in11(reg_weight16_32_1), .weight_in12(reg_weight16_32_2), .activation_in11(reg_activation17_31_1), .activation_in21(reg_activation17_31_2), .reg_partial_sum21(reg_psum17_32_1), .reg_partial_sum22(reg_psum17_32_2), .reg_weight21(reg_weight17_32_1), .reg_weight22(reg_weight17_32_2), .weight_en(weight_en));
SA22 U18_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_1_1), .partial_sum_in12(reg_psum17_1_2), .weight_in11(reg_weight17_1_1), .weight_in12(reg_weight17_1_2), .activation_in11(in_activation18_1_1), .activation_in21(in_activation18_1_2), .reg_partial_sum21(reg_psum18_1_1), .reg_partial_sum22(reg_psum18_1_2), .reg_weight21(reg_weight18_1_1), .reg_weight22(reg_weight18_1_2), .reg_activation12(reg_activation18_1_1), .reg_activation22(reg_activation18_1_2), .weight_en(weight_en));
SA22 U18_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_2_1), .partial_sum_in12(reg_psum17_2_2), .weight_in11(reg_weight17_2_1), .weight_in12(reg_weight17_2_2), .activation_in11(reg_activation18_1_1), .activation_in21(reg_activation18_1_2), .reg_partial_sum21(reg_psum18_2_1), .reg_partial_sum22(reg_psum18_2_2), .reg_weight21(reg_weight18_2_1), .reg_weight22(reg_weight18_2_2), .reg_activation12(reg_activation18_2_1), .reg_activation22(reg_activation18_2_2), .weight_en(weight_en));
SA22 U18_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_3_1), .partial_sum_in12(reg_psum17_3_2), .weight_in11(reg_weight17_3_1), .weight_in12(reg_weight17_3_2), .activation_in11(reg_activation18_2_1), .activation_in21(reg_activation18_2_2), .reg_partial_sum21(reg_psum18_3_1), .reg_partial_sum22(reg_psum18_3_2), .reg_weight21(reg_weight18_3_1), .reg_weight22(reg_weight18_3_2), .reg_activation12(reg_activation18_3_1), .reg_activation22(reg_activation18_3_2), .weight_en(weight_en));
SA22 U18_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_4_1), .partial_sum_in12(reg_psum17_4_2), .weight_in11(reg_weight17_4_1), .weight_in12(reg_weight17_4_2), .activation_in11(reg_activation18_3_1), .activation_in21(reg_activation18_3_2), .reg_partial_sum21(reg_psum18_4_1), .reg_partial_sum22(reg_psum18_4_2), .reg_weight21(reg_weight18_4_1), .reg_weight22(reg_weight18_4_2), .reg_activation12(reg_activation18_4_1), .reg_activation22(reg_activation18_4_2), .weight_en(weight_en));
SA22 U18_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_5_1), .partial_sum_in12(reg_psum17_5_2), .weight_in11(reg_weight17_5_1), .weight_in12(reg_weight17_5_2), .activation_in11(reg_activation18_4_1), .activation_in21(reg_activation18_4_2), .reg_partial_sum21(reg_psum18_5_1), .reg_partial_sum22(reg_psum18_5_2), .reg_weight21(reg_weight18_5_1), .reg_weight22(reg_weight18_5_2), .reg_activation12(reg_activation18_5_1), .reg_activation22(reg_activation18_5_2), .weight_en(weight_en));
SA22 U18_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_6_1), .partial_sum_in12(reg_psum17_6_2), .weight_in11(reg_weight17_6_1), .weight_in12(reg_weight17_6_2), .activation_in11(reg_activation18_5_1), .activation_in21(reg_activation18_5_2), .reg_partial_sum21(reg_psum18_6_1), .reg_partial_sum22(reg_psum18_6_2), .reg_weight21(reg_weight18_6_1), .reg_weight22(reg_weight18_6_2), .reg_activation12(reg_activation18_6_1), .reg_activation22(reg_activation18_6_2), .weight_en(weight_en));
SA22 U18_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_7_1), .partial_sum_in12(reg_psum17_7_2), .weight_in11(reg_weight17_7_1), .weight_in12(reg_weight17_7_2), .activation_in11(reg_activation18_6_1), .activation_in21(reg_activation18_6_2), .reg_partial_sum21(reg_psum18_7_1), .reg_partial_sum22(reg_psum18_7_2), .reg_weight21(reg_weight18_7_1), .reg_weight22(reg_weight18_7_2), .reg_activation12(reg_activation18_7_1), .reg_activation22(reg_activation18_7_2), .weight_en(weight_en));
SA22 U18_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_8_1), .partial_sum_in12(reg_psum17_8_2), .weight_in11(reg_weight17_8_1), .weight_in12(reg_weight17_8_2), .activation_in11(reg_activation18_7_1), .activation_in21(reg_activation18_7_2), .reg_partial_sum21(reg_psum18_8_1), .reg_partial_sum22(reg_psum18_8_2), .reg_weight21(reg_weight18_8_1), .reg_weight22(reg_weight18_8_2), .reg_activation12(reg_activation18_8_1), .reg_activation22(reg_activation18_8_2), .weight_en(weight_en));
SA22 U18_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_9_1), .partial_sum_in12(reg_psum17_9_2), .weight_in11(reg_weight17_9_1), .weight_in12(reg_weight17_9_2), .activation_in11(reg_activation18_8_1), .activation_in21(reg_activation18_8_2), .reg_partial_sum21(reg_psum18_9_1), .reg_partial_sum22(reg_psum18_9_2), .reg_weight21(reg_weight18_9_1), .reg_weight22(reg_weight18_9_2), .reg_activation12(reg_activation18_9_1), .reg_activation22(reg_activation18_9_2), .weight_en(weight_en));
SA22 U18_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_10_1), .partial_sum_in12(reg_psum17_10_2), .weight_in11(reg_weight17_10_1), .weight_in12(reg_weight17_10_2), .activation_in11(reg_activation18_9_1), .activation_in21(reg_activation18_9_2), .reg_partial_sum21(reg_psum18_10_1), .reg_partial_sum22(reg_psum18_10_2), .reg_weight21(reg_weight18_10_1), .reg_weight22(reg_weight18_10_2), .reg_activation12(reg_activation18_10_1), .reg_activation22(reg_activation18_10_2), .weight_en(weight_en));
SA22 U18_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_11_1), .partial_sum_in12(reg_psum17_11_2), .weight_in11(reg_weight17_11_1), .weight_in12(reg_weight17_11_2), .activation_in11(reg_activation18_10_1), .activation_in21(reg_activation18_10_2), .reg_partial_sum21(reg_psum18_11_1), .reg_partial_sum22(reg_psum18_11_2), .reg_weight21(reg_weight18_11_1), .reg_weight22(reg_weight18_11_2), .reg_activation12(reg_activation18_11_1), .reg_activation22(reg_activation18_11_2), .weight_en(weight_en));
SA22 U18_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_12_1), .partial_sum_in12(reg_psum17_12_2), .weight_in11(reg_weight17_12_1), .weight_in12(reg_weight17_12_2), .activation_in11(reg_activation18_11_1), .activation_in21(reg_activation18_11_2), .reg_partial_sum21(reg_psum18_12_1), .reg_partial_sum22(reg_psum18_12_2), .reg_weight21(reg_weight18_12_1), .reg_weight22(reg_weight18_12_2), .reg_activation12(reg_activation18_12_1), .reg_activation22(reg_activation18_12_2), .weight_en(weight_en));
SA22 U18_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_13_1), .partial_sum_in12(reg_psum17_13_2), .weight_in11(reg_weight17_13_1), .weight_in12(reg_weight17_13_2), .activation_in11(reg_activation18_12_1), .activation_in21(reg_activation18_12_2), .reg_partial_sum21(reg_psum18_13_1), .reg_partial_sum22(reg_psum18_13_2), .reg_weight21(reg_weight18_13_1), .reg_weight22(reg_weight18_13_2), .reg_activation12(reg_activation18_13_1), .reg_activation22(reg_activation18_13_2), .weight_en(weight_en));
SA22 U18_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_14_1), .partial_sum_in12(reg_psum17_14_2), .weight_in11(reg_weight17_14_1), .weight_in12(reg_weight17_14_2), .activation_in11(reg_activation18_13_1), .activation_in21(reg_activation18_13_2), .reg_partial_sum21(reg_psum18_14_1), .reg_partial_sum22(reg_psum18_14_2), .reg_weight21(reg_weight18_14_1), .reg_weight22(reg_weight18_14_2), .reg_activation12(reg_activation18_14_1), .reg_activation22(reg_activation18_14_2), .weight_en(weight_en));
SA22 U18_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_15_1), .partial_sum_in12(reg_psum17_15_2), .weight_in11(reg_weight17_15_1), .weight_in12(reg_weight17_15_2), .activation_in11(reg_activation18_14_1), .activation_in21(reg_activation18_14_2), .reg_partial_sum21(reg_psum18_15_1), .reg_partial_sum22(reg_psum18_15_2), .reg_weight21(reg_weight18_15_1), .reg_weight22(reg_weight18_15_2), .reg_activation12(reg_activation18_15_1), .reg_activation22(reg_activation18_15_2), .weight_en(weight_en));
SA22 U18_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_16_1), .partial_sum_in12(reg_psum17_16_2), .weight_in11(reg_weight17_16_1), .weight_in12(reg_weight17_16_2), .activation_in11(reg_activation18_15_1), .activation_in21(reg_activation18_15_2), .reg_partial_sum21(reg_psum18_16_1), .reg_partial_sum22(reg_psum18_16_2), .reg_weight21(reg_weight18_16_1), .reg_weight22(reg_weight18_16_2), .reg_activation12(reg_activation18_16_1), .reg_activation22(reg_activation18_16_2), .weight_en(weight_en));
SA22 U18_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_17_1), .partial_sum_in12(reg_psum17_17_2), .weight_in11(reg_weight17_17_1), .weight_in12(reg_weight17_17_2), .activation_in11(reg_activation18_16_1), .activation_in21(reg_activation18_16_2), .reg_partial_sum21(reg_psum18_17_1), .reg_partial_sum22(reg_psum18_17_2), .reg_weight21(reg_weight18_17_1), .reg_weight22(reg_weight18_17_2), .reg_activation12(reg_activation18_17_1), .reg_activation22(reg_activation18_17_2), .weight_en(weight_en));
SA22 U18_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_18_1), .partial_sum_in12(reg_psum17_18_2), .weight_in11(reg_weight17_18_1), .weight_in12(reg_weight17_18_2), .activation_in11(reg_activation18_17_1), .activation_in21(reg_activation18_17_2), .reg_partial_sum21(reg_psum18_18_1), .reg_partial_sum22(reg_psum18_18_2), .reg_weight21(reg_weight18_18_1), .reg_weight22(reg_weight18_18_2), .reg_activation12(reg_activation18_18_1), .reg_activation22(reg_activation18_18_2), .weight_en(weight_en));
SA22 U18_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_19_1), .partial_sum_in12(reg_psum17_19_2), .weight_in11(reg_weight17_19_1), .weight_in12(reg_weight17_19_2), .activation_in11(reg_activation18_18_1), .activation_in21(reg_activation18_18_2), .reg_partial_sum21(reg_psum18_19_1), .reg_partial_sum22(reg_psum18_19_2), .reg_weight21(reg_weight18_19_1), .reg_weight22(reg_weight18_19_2), .reg_activation12(reg_activation18_19_1), .reg_activation22(reg_activation18_19_2), .weight_en(weight_en));
SA22 U18_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_20_1), .partial_sum_in12(reg_psum17_20_2), .weight_in11(reg_weight17_20_1), .weight_in12(reg_weight17_20_2), .activation_in11(reg_activation18_19_1), .activation_in21(reg_activation18_19_2), .reg_partial_sum21(reg_psum18_20_1), .reg_partial_sum22(reg_psum18_20_2), .reg_weight21(reg_weight18_20_1), .reg_weight22(reg_weight18_20_2), .reg_activation12(reg_activation18_20_1), .reg_activation22(reg_activation18_20_2), .weight_en(weight_en));
SA22 U18_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_21_1), .partial_sum_in12(reg_psum17_21_2), .weight_in11(reg_weight17_21_1), .weight_in12(reg_weight17_21_2), .activation_in11(reg_activation18_20_1), .activation_in21(reg_activation18_20_2), .reg_partial_sum21(reg_psum18_21_1), .reg_partial_sum22(reg_psum18_21_2), .reg_weight21(reg_weight18_21_1), .reg_weight22(reg_weight18_21_2), .reg_activation12(reg_activation18_21_1), .reg_activation22(reg_activation18_21_2), .weight_en(weight_en));
SA22 U18_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_22_1), .partial_sum_in12(reg_psum17_22_2), .weight_in11(reg_weight17_22_1), .weight_in12(reg_weight17_22_2), .activation_in11(reg_activation18_21_1), .activation_in21(reg_activation18_21_2), .reg_partial_sum21(reg_psum18_22_1), .reg_partial_sum22(reg_psum18_22_2), .reg_weight21(reg_weight18_22_1), .reg_weight22(reg_weight18_22_2), .reg_activation12(reg_activation18_22_1), .reg_activation22(reg_activation18_22_2), .weight_en(weight_en));
SA22 U18_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_23_1), .partial_sum_in12(reg_psum17_23_2), .weight_in11(reg_weight17_23_1), .weight_in12(reg_weight17_23_2), .activation_in11(reg_activation18_22_1), .activation_in21(reg_activation18_22_2), .reg_partial_sum21(reg_psum18_23_1), .reg_partial_sum22(reg_psum18_23_2), .reg_weight21(reg_weight18_23_1), .reg_weight22(reg_weight18_23_2), .reg_activation12(reg_activation18_23_1), .reg_activation22(reg_activation18_23_2), .weight_en(weight_en));
SA22 U18_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_24_1), .partial_sum_in12(reg_psum17_24_2), .weight_in11(reg_weight17_24_1), .weight_in12(reg_weight17_24_2), .activation_in11(reg_activation18_23_1), .activation_in21(reg_activation18_23_2), .reg_partial_sum21(reg_psum18_24_1), .reg_partial_sum22(reg_psum18_24_2), .reg_weight21(reg_weight18_24_1), .reg_weight22(reg_weight18_24_2), .reg_activation12(reg_activation18_24_1), .reg_activation22(reg_activation18_24_2), .weight_en(weight_en));
SA22 U18_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_25_1), .partial_sum_in12(reg_psum17_25_2), .weight_in11(reg_weight17_25_1), .weight_in12(reg_weight17_25_2), .activation_in11(reg_activation18_24_1), .activation_in21(reg_activation18_24_2), .reg_partial_sum21(reg_psum18_25_1), .reg_partial_sum22(reg_psum18_25_2), .reg_weight21(reg_weight18_25_1), .reg_weight22(reg_weight18_25_2), .reg_activation12(reg_activation18_25_1), .reg_activation22(reg_activation18_25_2), .weight_en(weight_en));
SA22 U18_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_26_1), .partial_sum_in12(reg_psum17_26_2), .weight_in11(reg_weight17_26_1), .weight_in12(reg_weight17_26_2), .activation_in11(reg_activation18_25_1), .activation_in21(reg_activation18_25_2), .reg_partial_sum21(reg_psum18_26_1), .reg_partial_sum22(reg_psum18_26_2), .reg_weight21(reg_weight18_26_1), .reg_weight22(reg_weight18_26_2), .reg_activation12(reg_activation18_26_1), .reg_activation22(reg_activation18_26_2), .weight_en(weight_en));
SA22 U18_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_27_1), .partial_sum_in12(reg_psum17_27_2), .weight_in11(reg_weight17_27_1), .weight_in12(reg_weight17_27_2), .activation_in11(reg_activation18_26_1), .activation_in21(reg_activation18_26_2), .reg_partial_sum21(reg_psum18_27_1), .reg_partial_sum22(reg_psum18_27_2), .reg_weight21(reg_weight18_27_1), .reg_weight22(reg_weight18_27_2), .reg_activation12(reg_activation18_27_1), .reg_activation22(reg_activation18_27_2), .weight_en(weight_en));
SA22 U18_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_28_1), .partial_sum_in12(reg_psum17_28_2), .weight_in11(reg_weight17_28_1), .weight_in12(reg_weight17_28_2), .activation_in11(reg_activation18_27_1), .activation_in21(reg_activation18_27_2), .reg_partial_sum21(reg_psum18_28_1), .reg_partial_sum22(reg_psum18_28_2), .reg_weight21(reg_weight18_28_1), .reg_weight22(reg_weight18_28_2), .reg_activation12(reg_activation18_28_1), .reg_activation22(reg_activation18_28_2), .weight_en(weight_en));
SA22 U18_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_29_1), .partial_sum_in12(reg_psum17_29_2), .weight_in11(reg_weight17_29_1), .weight_in12(reg_weight17_29_2), .activation_in11(reg_activation18_28_1), .activation_in21(reg_activation18_28_2), .reg_partial_sum21(reg_psum18_29_1), .reg_partial_sum22(reg_psum18_29_2), .reg_weight21(reg_weight18_29_1), .reg_weight22(reg_weight18_29_2), .reg_activation12(reg_activation18_29_1), .reg_activation22(reg_activation18_29_2), .weight_en(weight_en));
SA22 U18_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_30_1), .partial_sum_in12(reg_psum17_30_2), .weight_in11(reg_weight17_30_1), .weight_in12(reg_weight17_30_2), .activation_in11(reg_activation18_29_1), .activation_in21(reg_activation18_29_2), .reg_partial_sum21(reg_psum18_30_1), .reg_partial_sum22(reg_psum18_30_2), .reg_weight21(reg_weight18_30_1), .reg_weight22(reg_weight18_30_2), .reg_activation12(reg_activation18_30_1), .reg_activation22(reg_activation18_30_2), .weight_en(weight_en));
SA22 U18_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_31_1), .partial_sum_in12(reg_psum17_31_2), .weight_in11(reg_weight17_31_1), .weight_in12(reg_weight17_31_2), .activation_in11(reg_activation18_30_1), .activation_in21(reg_activation18_30_2), .reg_partial_sum21(reg_psum18_31_1), .reg_partial_sum22(reg_psum18_31_2), .reg_weight21(reg_weight18_31_1), .reg_weight22(reg_weight18_31_2), .reg_activation12(reg_activation18_31_1), .reg_activation22(reg_activation18_31_2), .weight_en(weight_en));
SA22 U18_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum17_32_1), .partial_sum_in12(reg_psum17_32_2), .weight_in11(reg_weight17_32_1), .weight_in12(reg_weight17_32_2), .activation_in11(reg_activation18_31_1), .activation_in21(reg_activation18_31_2), .reg_partial_sum21(reg_psum18_32_1), .reg_partial_sum22(reg_psum18_32_2), .reg_weight21(reg_weight18_32_1), .reg_weight22(reg_weight18_32_2), .weight_en(weight_en));
SA22 U19_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_1_1), .partial_sum_in12(reg_psum18_1_2), .weight_in11(reg_weight18_1_1), .weight_in12(reg_weight18_1_2), .activation_in11(in_activation19_1_1), .activation_in21(in_activation19_1_2), .reg_partial_sum21(reg_psum19_1_1), .reg_partial_sum22(reg_psum19_1_2), .reg_weight21(reg_weight19_1_1), .reg_weight22(reg_weight19_1_2), .reg_activation12(reg_activation19_1_1), .reg_activation22(reg_activation19_1_2), .weight_en(weight_en));
SA22 U19_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_2_1), .partial_sum_in12(reg_psum18_2_2), .weight_in11(reg_weight18_2_1), .weight_in12(reg_weight18_2_2), .activation_in11(reg_activation19_1_1), .activation_in21(reg_activation19_1_2), .reg_partial_sum21(reg_psum19_2_1), .reg_partial_sum22(reg_psum19_2_2), .reg_weight21(reg_weight19_2_1), .reg_weight22(reg_weight19_2_2), .reg_activation12(reg_activation19_2_1), .reg_activation22(reg_activation19_2_2), .weight_en(weight_en));
SA22 U19_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_3_1), .partial_sum_in12(reg_psum18_3_2), .weight_in11(reg_weight18_3_1), .weight_in12(reg_weight18_3_2), .activation_in11(reg_activation19_2_1), .activation_in21(reg_activation19_2_2), .reg_partial_sum21(reg_psum19_3_1), .reg_partial_sum22(reg_psum19_3_2), .reg_weight21(reg_weight19_3_1), .reg_weight22(reg_weight19_3_2), .reg_activation12(reg_activation19_3_1), .reg_activation22(reg_activation19_3_2), .weight_en(weight_en));
SA22 U19_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_4_1), .partial_sum_in12(reg_psum18_4_2), .weight_in11(reg_weight18_4_1), .weight_in12(reg_weight18_4_2), .activation_in11(reg_activation19_3_1), .activation_in21(reg_activation19_3_2), .reg_partial_sum21(reg_psum19_4_1), .reg_partial_sum22(reg_psum19_4_2), .reg_weight21(reg_weight19_4_1), .reg_weight22(reg_weight19_4_2), .reg_activation12(reg_activation19_4_1), .reg_activation22(reg_activation19_4_2), .weight_en(weight_en));
SA22 U19_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_5_1), .partial_sum_in12(reg_psum18_5_2), .weight_in11(reg_weight18_5_1), .weight_in12(reg_weight18_5_2), .activation_in11(reg_activation19_4_1), .activation_in21(reg_activation19_4_2), .reg_partial_sum21(reg_psum19_5_1), .reg_partial_sum22(reg_psum19_5_2), .reg_weight21(reg_weight19_5_1), .reg_weight22(reg_weight19_5_2), .reg_activation12(reg_activation19_5_1), .reg_activation22(reg_activation19_5_2), .weight_en(weight_en));
SA22 U19_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_6_1), .partial_sum_in12(reg_psum18_6_2), .weight_in11(reg_weight18_6_1), .weight_in12(reg_weight18_6_2), .activation_in11(reg_activation19_5_1), .activation_in21(reg_activation19_5_2), .reg_partial_sum21(reg_psum19_6_1), .reg_partial_sum22(reg_psum19_6_2), .reg_weight21(reg_weight19_6_1), .reg_weight22(reg_weight19_6_2), .reg_activation12(reg_activation19_6_1), .reg_activation22(reg_activation19_6_2), .weight_en(weight_en));
SA22 U19_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_7_1), .partial_sum_in12(reg_psum18_7_2), .weight_in11(reg_weight18_7_1), .weight_in12(reg_weight18_7_2), .activation_in11(reg_activation19_6_1), .activation_in21(reg_activation19_6_2), .reg_partial_sum21(reg_psum19_7_1), .reg_partial_sum22(reg_psum19_7_2), .reg_weight21(reg_weight19_7_1), .reg_weight22(reg_weight19_7_2), .reg_activation12(reg_activation19_7_1), .reg_activation22(reg_activation19_7_2), .weight_en(weight_en));
SA22 U19_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_8_1), .partial_sum_in12(reg_psum18_8_2), .weight_in11(reg_weight18_8_1), .weight_in12(reg_weight18_8_2), .activation_in11(reg_activation19_7_1), .activation_in21(reg_activation19_7_2), .reg_partial_sum21(reg_psum19_8_1), .reg_partial_sum22(reg_psum19_8_2), .reg_weight21(reg_weight19_8_1), .reg_weight22(reg_weight19_8_2), .reg_activation12(reg_activation19_8_1), .reg_activation22(reg_activation19_8_2), .weight_en(weight_en));
SA22 U19_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_9_1), .partial_sum_in12(reg_psum18_9_2), .weight_in11(reg_weight18_9_1), .weight_in12(reg_weight18_9_2), .activation_in11(reg_activation19_8_1), .activation_in21(reg_activation19_8_2), .reg_partial_sum21(reg_psum19_9_1), .reg_partial_sum22(reg_psum19_9_2), .reg_weight21(reg_weight19_9_1), .reg_weight22(reg_weight19_9_2), .reg_activation12(reg_activation19_9_1), .reg_activation22(reg_activation19_9_2), .weight_en(weight_en));
SA22 U19_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_10_1), .partial_sum_in12(reg_psum18_10_2), .weight_in11(reg_weight18_10_1), .weight_in12(reg_weight18_10_2), .activation_in11(reg_activation19_9_1), .activation_in21(reg_activation19_9_2), .reg_partial_sum21(reg_psum19_10_1), .reg_partial_sum22(reg_psum19_10_2), .reg_weight21(reg_weight19_10_1), .reg_weight22(reg_weight19_10_2), .reg_activation12(reg_activation19_10_1), .reg_activation22(reg_activation19_10_2), .weight_en(weight_en));
SA22 U19_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_11_1), .partial_sum_in12(reg_psum18_11_2), .weight_in11(reg_weight18_11_1), .weight_in12(reg_weight18_11_2), .activation_in11(reg_activation19_10_1), .activation_in21(reg_activation19_10_2), .reg_partial_sum21(reg_psum19_11_1), .reg_partial_sum22(reg_psum19_11_2), .reg_weight21(reg_weight19_11_1), .reg_weight22(reg_weight19_11_2), .reg_activation12(reg_activation19_11_1), .reg_activation22(reg_activation19_11_2), .weight_en(weight_en));
SA22 U19_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_12_1), .partial_sum_in12(reg_psum18_12_2), .weight_in11(reg_weight18_12_1), .weight_in12(reg_weight18_12_2), .activation_in11(reg_activation19_11_1), .activation_in21(reg_activation19_11_2), .reg_partial_sum21(reg_psum19_12_1), .reg_partial_sum22(reg_psum19_12_2), .reg_weight21(reg_weight19_12_1), .reg_weight22(reg_weight19_12_2), .reg_activation12(reg_activation19_12_1), .reg_activation22(reg_activation19_12_2), .weight_en(weight_en));
SA22 U19_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_13_1), .partial_sum_in12(reg_psum18_13_2), .weight_in11(reg_weight18_13_1), .weight_in12(reg_weight18_13_2), .activation_in11(reg_activation19_12_1), .activation_in21(reg_activation19_12_2), .reg_partial_sum21(reg_psum19_13_1), .reg_partial_sum22(reg_psum19_13_2), .reg_weight21(reg_weight19_13_1), .reg_weight22(reg_weight19_13_2), .reg_activation12(reg_activation19_13_1), .reg_activation22(reg_activation19_13_2), .weight_en(weight_en));
SA22 U19_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_14_1), .partial_sum_in12(reg_psum18_14_2), .weight_in11(reg_weight18_14_1), .weight_in12(reg_weight18_14_2), .activation_in11(reg_activation19_13_1), .activation_in21(reg_activation19_13_2), .reg_partial_sum21(reg_psum19_14_1), .reg_partial_sum22(reg_psum19_14_2), .reg_weight21(reg_weight19_14_1), .reg_weight22(reg_weight19_14_2), .reg_activation12(reg_activation19_14_1), .reg_activation22(reg_activation19_14_2), .weight_en(weight_en));
SA22 U19_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_15_1), .partial_sum_in12(reg_psum18_15_2), .weight_in11(reg_weight18_15_1), .weight_in12(reg_weight18_15_2), .activation_in11(reg_activation19_14_1), .activation_in21(reg_activation19_14_2), .reg_partial_sum21(reg_psum19_15_1), .reg_partial_sum22(reg_psum19_15_2), .reg_weight21(reg_weight19_15_1), .reg_weight22(reg_weight19_15_2), .reg_activation12(reg_activation19_15_1), .reg_activation22(reg_activation19_15_2), .weight_en(weight_en));
SA22 U19_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_16_1), .partial_sum_in12(reg_psum18_16_2), .weight_in11(reg_weight18_16_1), .weight_in12(reg_weight18_16_2), .activation_in11(reg_activation19_15_1), .activation_in21(reg_activation19_15_2), .reg_partial_sum21(reg_psum19_16_1), .reg_partial_sum22(reg_psum19_16_2), .reg_weight21(reg_weight19_16_1), .reg_weight22(reg_weight19_16_2), .reg_activation12(reg_activation19_16_1), .reg_activation22(reg_activation19_16_2), .weight_en(weight_en));
SA22 U19_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_17_1), .partial_sum_in12(reg_psum18_17_2), .weight_in11(reg_weight18_17_1), .weight_in12(reg_weight18_17_2), .activation_in11(reg_activation19_16_1), .activation_in21(reg_activation19_16_2), .reg_partial_sum21(reg_psum19_17_1), .reg_partial_sum22(reg_psum19_17_2), .reg_weight21(reg_weight19_17_1), .reg_weight22(reg_weight19_17_2), .reg_activation12(reg_activation19_17_1), .reg_activation22(reg_activation19_17_2), .weight_en(weight_en));
SA22 U19_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_18_1), .partial_sum_in12(reg_psum18_18_2), .weight_in11(reg_weight18_18_1), .weight_in12(reg_weight18_18_2), .activation_in11(reg_activation19_17_1), .activation_in21(reg_activation19_17_2), .reg_partial_sum21(reg_psum19_18_1), .reg_partial_sum22(reg_psum19_18_2), .reg_weight21(reg_weight19_18_1), .reg_weight22(reg_weight19_18_2), .reg_activation12(reg_activation19_18_1), .reg_activation22(reg_activation19_18_2), .weight_en(weight_en));
SA22 U19_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_19_1), .partial_sum_in12(reg_psum18_19_2), .weight_in11(reg_weight18_19_1), .weight_in12(reg_weight18_19_2), .activation_in11(reg_activation19_18_1), .activation_in21(reg_activation19_18_2), .reg_partial_sum21(reg_psum19_19_1), .reg_partial_sum22(reg_psum19_19_2), .reg_weight21(reg_weight19_19_1), .reg_weight22(reg_weight19_19_2), .reg_activation12(reg_activation19_19_1), .reg_activation22(reg_activation19_19_2), .weight_en(weight_en));
SA22 U19_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_20_1), .partial_sum_in12(reg_psum18_20_2), .weight_in11(reg_weight18_20_1), .weight_in12(reg_weight18_20_2), .activation_in11(reg_activation19_19_1), .activation_in21(reg_activation19_19_2), .reg_partial_sum21(reg_psum19_20_1), .reg_partial_sum22(reg_psum19_20_2), .reg_weight21(reg_weight19_20_1), .reg_weight22(reg_weight19_20_2), .reg_activation12(reg_activation19_20_1), .reg_activation22(reg_activation19_20_2), .weight_en(weight_en));
SA22 U19_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_21_1), .partial_sum_in12(reg_psum18_21_2), .weight_in11(reg_weight18_21_1), .weight_in12(reg_weight18_21_2), .activation_in11(reg_activation19_20_1), .activation_in21(reg_activation19_20_2), .reg_partial_sum21(reg_psum19_21_1), .reg_partial_sum22(reg_psum19_21_2), .reg_weight21(reg_weight19_21_1), .reg_weight22(reg_weight19_21_2), .reg_activation12(reg_activation19_21_1), .reg_activation22(reg_activation19_21_2), .weight_en(weight_en));
SA22 U19_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_22_1), .partial_sum_in12(reg_psum18_22_2), .weight_in11(reg_weight18_22_1), .weight_in12(reg_weight18_22_2), .activation_in11(reg_activation19_21_1), .activation_in21(reg_activation19_21_2), .reg_partial_sum21(reg_psum19_22_1), .reg_partial_sum22(reg_psum19_22_2), .reg_weight21(reg_weight19_22_1), .reg_weight22(reg_weight19_22_2), .reg_activation12(reg_activation19_22_1), .reg_activation22(reg_activation19_22_2), .weight_en(weight_en));
SA22 U19_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_23_1), .partial_sum_in12(reg_psum18_23_2), .weight_in11(reg_weight18_23_1), .weight_in12(reg_weight18_23_2), .activation_in11(reg_activation19_22_1), .activation_in21(reg_activation19_22_2), .reg_partial_sum21(reg_psum19_23_1), .reg_partial_sum22(reg_psum19_23_2), .reg_weight21(reg_weight19_23_1), .reg_weight22(reg_weight19_23_2), .reg_activation12(reg_activation19_23_1), .reg_activation22(reg_activation19_23_2), .weight_en(weight_en));
SA22 U19_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_24_1), .partial_sum_in12(reg_psum18_24_2), .weight_in11(reg_weight18_24_1), .weight_in12(reg_weight18_24_2), .activation_in11(reg_activation19_23_1), .activation_in21(reg_activation19_23_2), .reg_partial_sum21(reg_psum19_24_1), .reg_partial_sum22(reg_psum19_24_2), .reg_weight21(reg_weight19_24_1), .reg_weight22(reg_weight19_24_2), .reg_activation12(reg_activation19_24_1), .reg_activation22(reg_activation19_24_2), .weight_en(weight_en));
SA22 U19_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_25_1), .partial_sum_in12(reg_psum18_25_2), .weight_in11(reg_weight18_25_1), .weight_in12(reg_weight18_25_2), .activation_in11(reg_activation19_24_1), .activation_in21(reg_activation19_24_2), .reg_partial_sum21(reg_psum19_25_1), .reg_partial_sum22(reg_psum19_25_2), .reg_weight21(reg_weight19_25_1), .reg_weight22(reg_weight19_25_2), .reg_activation12(reg_activation19_25_1), .reg_activation22(reg_activation19_25_2), .weight_en(weight_en));
SA22 U19_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_26_1), .partial_sum_in12(reg_psum18_26_2), .weight_in11(reg_weight18_26_1), .weight_in12(reg_weight18_26_2), .activation_in11(reg_activation19_25_1), .activation_in21(reg_activation19_25_2), .reg_partial_sum21(reg_psum19_26_1), .reg_partial_sum22(reg_psum19_26_2), .reg_weight21(reg_weight19_26_1), .reg_weight22(reg_weight19_26_2), .reg_activation12(reg_activation19_26_1), .reg_activation22(reg_activation19_26_2), .weight_en(weight_en));
SA22 U19_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_27_1), .partial_sum_in12(reg_psum18_27_2), .weight_in11(reg_weight18_27_1), .weight_in12(reg_weight18_27_2), .activation_in11(reg_activation19_26_1), .activation_in21(reg_activation19_26_2), .reg_partial_sum21(reg_psum19_27_1), .reg_partial_sum22(reg_psum19_27_2), .reg_weight21(reg_weight19_27_1), .reg_weight22(reg_weight19_27_2), .reg_activation12(reg_activation19_27_1), .reg_activation22(reg_activation19_27_2), .weight_en(weight_en));
SA22 U19_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_28_1), .partial_sum_in12(reg_psum18_28_2), .weight_in11(reg_weight18_28_1), .weight_in12(reg_weight18_28_2), .activation_in11(reg_activation19_27_1), .activation_in21(reg_activation19_27_2), .reg_partial_sum21(reg_psum19_28_1), .reg_partial_sum22(reg_psum19_28_2), .reg_weight21(reg_weight19_28_1), .reg_weight22(reg_weight19_28_2), .reg_activation12(reg_activation19_28_1), .reg_activation22(reg_activation19_28_2), .weight_en(weight_en));
SA22 U19_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_29_1), .partial_sum_in12(reg_psum18_29_2), .weight_in11(reg_weight18_29_1), .weight_in12(reg_weight18_29_2), .activation_in11(reg_activation19_28_1), .activation_in21(reg_activation19_28_2), .reg_partial_sum21(reg_psum19_29_1), .reg_partial_sum22(reg_psum19_29_2), .reg_weight21(reg_weight19_29_1), .reg_weight22(reg_weight19_29_2), .reg_activation12(reg_activation19_29_1), .reg_activation22(reg_activation19_29_2), .weight_en(weight_en));
SA22 U19_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_30_1), .partial_sum_in12(reg_psum18_30_2), .weight_in11(reg_weight18_30_1), .weight_in12(reg_weight18_30_2), .activation_in11(reg_activation19_29_1), .activation_in21(reg_activation19_29_2), .reg_partial_sum21(reg_psum19_30_1), .reg_partial_sum22(reg_psum19_30_2), .reg_weight21(reg_weight19_30_1), .reg_weight22(reg_weight19_30_2), .reg_activation12(reg_activation19_30_1), .reg_activation22(reg_activation19_30_2), .weight_en(weight_en));
SA22 U19_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_31_1), .partial_sum_in12(reg_psum18_31_2), .weight_in11(reg_weight18_31_1), .weight_in12(reg_weight18_31_2), .activation_in11(reg_activation19_30_1), .activation_in21(reg_activation19_30_2), .reg_partial_sum21(reg_psum19_31_1), .reg_partial_sum22(reg_psum19_31_2), .reg_weight21(reg_weight19_31_1), .reg_weight22(reg_weight19_31_2), .reg_activation12(reg_activation19_31_1), .reg_activation22(reg_activation19_31_2), .weight_en(weight_en));
SA22 U19_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum18_32_1), .partial_sum_in12(reg_psum18_32_2), .weight_in11(reg_weight18_32_1), .weight_in12(reg_weight18_32_2), .activation_in11(reg_activation19_31_1), .activation_in21(reg_activation19_31_2), .reg_partial_sum21(reg_psum19_32_1), .reg_partial_sum22(reg_psum19_32_2), .reg_weight21(reg_weight19_32_1), .reg_weight22(reg_weight19_32_2), .weight_en(weight_en));
SA22 U20_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_1_1), .partial_sum_in12(reg_psum19_1_2), .weight_in11(reg_weight19_1_1), .weight_in12(reg_weight19_1_2), .activation_in11(in_activation20_1_1), .activation_in21(in_activation20_1_2), .reg_partial_sum21(reg_psum20_1_1), .reg_partial_sum22(reg_psum20_1_2), .reg_weight21(reg_weight20_1_1), .reg_weight22(reg_weight20_1_2), .reg_activation12(reg_activation20_1_1), .reg_activation22(reg_activation20_1_2), .weight_en(weight_en));
SA22 U20_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_2_1), .partial_sum_in12(reg_psum19_2_2), .weight_in11(reg_weight19_2_1), .weight_in12(reg_weight19_2_2), .activation_in11(reg_activation20_1_1), .activation_in21(reg_activation20_1_2), .reg_partial_sum21(reg_psum20_2_1), .reg_partial_sum22(reg_psum20_2_2), .reg_weight21(reg_weight20_2_1), .reg_weight22(reg_weight20_2_2), .reg_activation12(reg_activation20_2_1), .reg_activation22(reg_activation20_2_2), .weight_en(weight_en));
SA22 U20_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_3_1), .partial_sum_in12(reg_psum19_3_2), .weight_in11(reg_weight19_3_1), .weight_in12(reg_weight19_3_2), .activation_in11(reg_activation20_2_1), .activation_in21(reg_activation20_2_2), .reg_partial_sum21(reg_psum20_3_1), .reg_partial_sum22(reg_psum20_3_2), .reg_weight21(reg_weight20_3_1), .reg_weight22(reg_weight20_3_2), .reg_activation12(reg_activation20_3_1), .reg_activation22(reg_activation20_3_2), .weight_en(weight_en));
SA22 U20_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_4_1), .partial_sum_in12(reg_psum19_4_2), .weight_in11(reg_weight19_4_1), .weight_in12(reg_weight19_4_2), .activation_in11(reg_activation20_3_1), .activation_in21(reg_activation20_3_2), .reg_partial_sum21(reg_psum20_4_1), .reg_partial_sum22(reg_psum20_4_2), .reg_weight21(reg_weight20_4_1), .reg_weight22(reg_weight20_4_2), .reg_activation12(reg_activation20_4_1), .reg_activation22(reg_activation20_4_2), .weight_en(weight_en));
SA22 U20_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_5_1), .partial_sum_in12(reg_psum19_5_2), .weight_in11(reg_weight19_5_1), .weight_in12(reg_weight19_5_2), .activation_in11(reg_activation20_4_1), .activation_in21(reg_activation20_4_2), .reg_partial_sum21(reg_psum20_5_1), .reg_partial_sum22(reg_psum20_5_2), .reg_weight21(reg_weight20_5_1), .reg_weight22(reg_weight20_5_2), .reg_activation12(reg_activation20_5_1), .reg_activation22(reg_activation20_5_2), .weight_en(weight_en));
SA22 U20_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_6_1), .partial_sum_in12(reg_psum19_6_2), .weight_in11(reg_weight19_6_1), .weight_in12(reg_weight19_6_2), .activation_in11(reg_activation20_5_1), .activation_in21(reg_activation20_5_2), .reg_partial_sum21(reg_psum20_6_1), .reg_partial_sum22(reg_psum20_6_2), .reg_weight21(reg_weight20_6_1), .reg_weight22(reg_weight20_6_2), .reg_activation12(reg_activation20_6_1), .reg_activation22(reg_activation20_6_2), .weight_en(weight_en));
SA22 U20_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_7_1), .partial_sum_in12(reg_psum19_7_2), .weight_in11(reg_weight19_7_1), .weight_in12(reg_weight19_7_2), .activation_in11(reg_activation20_6_1), .activation_in21(reg_activation20_6_2), .reg_partial_sum21(reg_psum20_7_1), .reg_partial_sum22(reg_psum20_7_2), .reg_weight21(reg_weight20_7_1), .reg_weight22(reg_weight20_7_2), .reg_activation12(reg_activation20_7_1), .reg_activation22(reg_activation20_7_2), .weight_en(weight_en));
SA22 U20_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_8_1), .partial_sum_in12(reg_psum19_8_2), .weight_in11(reg_weight19_8_1), .weight_in12(reg_weight19_8_2), .activation_in11(reg_activation20_7_1), .activation_in21(reg_activation20_7_2), .reg_partial_sum21(reg_psum20_8_1), .reg_partial_sum22(reg_psum20_8_2), .reg_weight21(reg_weight20_8_1), .reg_weight22(reg_weight20_8_2), .reg_activation12(reg_activation20_8_1), .reg_activation22(reg_activation20_8_2), .weight_en(weight_en));
SA22 U20_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_9_1), .partial_sum_in12(reg_psum19_9_2), .weight_in11(reg_weight19_9_1), .weight_in12(reg_weight19_9_2), .activation_in11(reg_activation20_8_1), .activation_in21(reg_activation20_8_2), .reg_partial_sum21(reg_psum20_9_1), .reg_partial_sum22(reg_psum20_9_2), .reg_weight21(reg_weight20_9_1), .reg_weight22(reg_weight20_9_2), .reg_activation12(reg_activation20_9_1), .reg_activation22(reg_activation20_9_2), .weight_en(weight_en));
SA22 U20_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_10_1), .partial_sum_in12(reg_psum19_10_2), .weight_in11(reg_weight19_10_1), .weight_in12(reg_weight19_10_2), .activation_in11(reg_activation20_9_1), .activation_in21(reg_activation20_9_2), .reg_partial_sum21(reg_psum20_10_1), .reg_partial_sum22(reg_psum20_10_2), .reg_weight21(reg_weight20_10_1), .reg_weight22(reg_weight20_10_2), .reg_activation12(reg_activation20_10_1), .reg_activation22(reg_activation20_10_2), .weight_en(weight_en));
SA22 U20_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_11_1), .partial_sum_in12(reg_psum19_11_2), .weight_in11(reg_weight19_11_1), .weight_in12(reg_weight19_11_2), .activation_in11(reg_activation20_10_1), .activation_in21(reg_activation20_10_2), .reg_partial_sum21(reg_psum20_11_1), .reg_partial_sum22(reg_psum20_11_2), .reg_weight21(reg_weight20_11_1), .reg_weight22(reg_weight20_11_2), .reg_activation12(reg_activation20_11_1), .reg_activation22(reg_activation20_11_2), .weight_en(weight_en));
SA22 U20_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_12_1), .partial_sum_in12(reg_psum19_12_2), .weight_in11(reg_weight19_12_1), .weight_in12(reg_weight19_12_2), .activation_in11(reg_activation20_11_1), .activation_in21(reg_activation20_11_2), .reg_partial_sum21(reg_psum20_12_1), .reg_partial_sum22(reg_psum20_12_2), .reg_weight21(reg_weight20_12_1), .reg_weight22(reg_weight20_12_2), .reg_activation12(reg_activation20_12_1), .reg_activation22(reg_activation20_12_2), .weight_en(weight_en));
SA22 U20_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_13_1), .partial_sum_in12(reg_psum19_13_2), .weight_in11(reg_weight19_13_1), .weight_in12(reg_weight19_13_2), .activation_in11(reg_activation20_12_1), .activation_in21(reg_activation20_12_2), .reg_partial_sum21(reg_psum20_13_1), .reg_partial_sum22(reg_psum20_13_2), .reg_weight21(reg_weight20_13_1), .reg_weight22(reg_weight20_13_2), .reg_activation12(reg_activation20_13_1), .reg_activation22(reg_activation20_13_2), .weight_en(weight_en));
SA22 U20_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_14_1), .partial_sum_in12(reg_psum19_14_2), .weight_in11(reg_weight19_14_1), .weight_in12(reg_weight19_14_2), .activation_in11(reg_activation20_13_1), .activation_in21(reg_activation20_13_2), .reg_partial_sum21(reg_psum20_14_1), .reg_partial_sum22(reg_psum20_14_2), .reg_weight21(reg_weight20_14_1), .reg_weight22(reg_weight20_14_2), .reg_activation12(reg_activation20_14_1), .reg_activation22(reg_activation20_14_2), .weight_en(weight_en));
SA22 U20_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_15_1), .partial_sum_in12(reg_psum19_15_2), .weight_in11(reg_weight19_15_1), .weight_in12(reg_weight19_15_2), .activation_in11(reg_activation20_14_1), .activation_in21(reg_activation20_14_2), .reg_partial_sum21(reg_psum20_15_1), .reg_partial_sum22(reg_psum20_15_2), .reg_weight21(reg_weight20_15_1), .reg_weight22(reg_weight20_15_2), .reg_activation12(reg_activation20_15_1), .reg_activation22(reg_activation20_15_2), .weight_en(weight_en));
SA22 U20_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_16_1), .partial_sum_in12(reg_psum19_16_2), .weight_in11(reg_weight19_16_1), .weight_in12(reg_weight19_16_2), .activation_in11(reg_activation20_15_1), .activation_in21(reg_activation20_15_2), .reg_partial_sum21(reg_psum20_16_1), .reg_partial_sum22(reg_psum20_16_2), .reg_weight21(reg_weight20_16_1), .reg_weight22(reg_weight20_16_2), .reg_activation12(reg_activation20_16_1), .reg_activation22(reg_activation20_16_2), .weight_en(weight_en));
SA22 U20_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_17_1), .partial_sum_in12(reg_psum19_17_2), .weight_in11(reg_weight19_17_1), .weight_in12(reg_weight19_17_2), .activation_in11(reg_activation20_16_1), .activation_in21(reg_activation20_16_2), .reg_partial_sum21(reg_psum20_17_1), .reg_partial_sum22(reg_psum20_17_2), .reg_weight21(reg_weight20_17_1), .reg_weight22(reg_weight20_17_2), .reg_activation12(reg_activation20_17_1), .reg_activation22(reg_activation20_17_2), .weight_en(weight_en));
SA22 U20_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_18_1), .partial_sum_in12(reg_psum19_18_2), .weight_in11(reg_weight19_18_1), .weight_in12(reg_weight19_18_2), .activation_in11(reg_activation20_17_1), .activation_in21(reg_activation20_17_2), .reg_partial_sum21(reg_psum20_18_1), .reg_partial_sum22(reg_psum20_18_2), .reg_weight21(reg_weight20_18_1), .reg_weight22(reg_weight20_18_2), .reg_activation12(reg_activation20_18_1), .reg_activation22(reg_activation20_18_2), .weight_en(weight_en));
SA22 U20_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_19_1), .partial_sum_in12(reg_psum19_19_2), .weight_in11(reg_weight19_19_1), .weight_in12(reg_weight19_19_2), .activation_in11(reg_activation20_18_1), .activation_in21(reg_activation20_18_2), .reg_partial_sum21(reg_psum20_19_1), .reg_partial_sum22(reg_psum20_19_2), .reg_weight21(reg_weight20_19_1), .reg_weight22(reg_weight20_19_2), .reg_activation12(reg_activation20_19_1), .reg_activation22(reg_activation20_19_2), .weight_en(weight_en));
SA22 U20_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_20_1), .partial_sum_in12(reg_psum19_20_2), .weight_in11(reg_weight19_20_1), .weight_in12(reg_weight19_20_2), .activation_in11(reg_activation20_19_1), .activation_in21(reg_activation20_19_2), .reg_partial_sum21(reg_psum20_20_1), .reg_partial_sum22(reg_psum20_20_2), .reg_weight21(reg_weight20_20_1), .reg_weight22(reg_weight20_20_2), .reg_activation12(reg_activation20_20_1), .reg_activation22(reg_activation20_20_2), .weight_en(weight_en));
SA22 U20_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_21_1), .partial_sum_in12(reg_psum19_21_2), .weight_in11(reg_weight19_21_1), .weight_in12(reg_weight19_21_2), .activation_in11(reg_activation20_20_1), .activation_in21(reg_activation20_20_2), .reg_partial_sum21(reg_psum20_21_1), .reg_partial_sum22(reg_psum20_21_2), .reg_weight21(reg_weight20_21_1), .reg_weight22(reg_weight20_21_2), .reg_activation12(reg_activation20_21_1), .reg_activation22(reg_activation20_21_2), .weight_en(weight_en));
SA22 U20_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_22_1), .partial_sum_in12(reg_psum19_22_2), .weight_in11(reg_weight19_22_1), .weight_in12(reg_weight19_22_2), .activation_in11(reg_activation20_21_1), .activation_in21(reg_activation20_21_2), .reg_partial_sum21(reg_psum20_22_1), .reg_partial_sum22(reg_psum20_22_2), .reg_weight21(reg_weight20_22_1), .reg_weight22(reg_weight20_22_2), .reg_activation12(reg_activation20_22_1), .reg_activation22(reg_activation20_22_2), .weight_en(weight_en));
SA22 U20_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_23_1), .partial_sum_in12(reg_psum19_23_2), .weight_in11(reg_weight19_23_1), .weight_in12(reg_weight19_23_2), .activation_in11(reg_activation20_22_1), .activation_in21(reg_activation20_22_2), .reg_partial_sum21(reg_psum20_23_1), .reg_partial_sum22(reg_psum20_23_2), .reg_weight21(reg_weight20_23_1), .reg_weight22(reg_weight20_23_2), .reg_activation12(reg_activation20_23_1), .reg_activation22(reg_activation20_23_2), .weight_en(weight_en));
SA22 U20_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_24_1), .partial_sum_in12(reg_psum19_24_2), .weight_in11(reg_weight19_24_1), .weight_in12(reg_weight19_24_2), .activation_in11(reg_activation20_23_1), .activation_in21(reg_activation20_23_2), .reg_partial_sum21(reg_psum20_24_1), .reg_partial_sum22(reg_psum20_24_2), .reg_weight21(reg_weight20_24_1), .reg_weight22(reg_weight20_24_2), .reg_activation12(reg_activation20_24_1), .reg_activation22(reg_activation20_24_2), .weight_en(weight_en));
SA22 U20_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_25_1), .partial_sum_in12(reg_psum19_25_2), .weight_in11(reg_weight19_25_1), .weight_in12(reg_weight19_25_2), .activation_in11(reg_activation20_24_1), .activation_in21(reg_activation20_24_2), .reg_partial_sum21(reg_psum20_25_1), .reg_partial_sum22(reg_psum20_25_2), .reg_weight21(reg_weight20_25_1), .reg_weight22(reg_weight20_25_2), .reg_activation12(reg_activation20_25_1), .reg_activation22(reg_activation20_25_2), .weight_en(weight_en));
SA22 U20_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_26_1), .partial_sum_in12(reg_psum19_26_2), .weight_in11(reg_weight19_26_1), .weight_in12(reg_weight19_26_2), .activation_in11(reg_activation20_25_1), .activation_in21(reg_activation20_25_2), .reg_partial_sum21(reg_psum20_26_1), .reg_partial_sum22(reg_psum20_26_2), .reg_weight21(reg_weight20_26_1), .reg_weight22(reg_weight20_26_2), .reg_activation12(reg_activation20_26_1), .reg_activation22(reg_activation20_26_2), .weight_en(weight_en));
SA22 U20_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_27_1), .partial_sum_in12(reg_psum19_27_2), .weight_in11(reg_weight19_27_1), .weight_in12(reg_weight19_27_2), .activation_in11(reg_activation20_26_1), .activation_in21(reg_activation20_26_2), .reg_partial_sum21(reg_psum20_27_1), .reg_partial_sum22(reg_psum20_27_2), .reg_weight21(reg_weight20_27_1), .reg_weight22(reg_weight20_27_2), .reg_activation12(reg_activation20_27_1), .reg_activation22(reg_activation20_27_2), .weight_en(weight_en));
SA22 U20_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_28_1), .partial_sum_in12(reg_psum19_28_2), .weight_in11(reg_weight19_28_1), .weight_in12(reg_weight19_28_2), .activation_in11(reg_activation20_27_1), .activation_in21(reg_activation20_27_2), .reg_partial_sum21(reg_psum20_28_1), .reg_partial_sum22(reg_psum20_28_2), .reg_weight21(reg_weight20_28_1), .reg_weight22(reg_weight20_28_2), .reg_activation12(reg_activation20_28_1), .reg_activation22(reg_activation20_28_2), .weight_en(weight_en));
SA22 U20_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_29_1), .partial_sum_in12(reg_psum19_29_2), .weight_in11(reg_weight19_29_1), .weight_in12(reg_weight19_29_2), .activation_in11(reg_activation20_28_1), .activation_in21(reg_activation20_28_2), .reg_partial_sum21(reg_psum20_29_1), .reg_partial_sum22(reg_psum20_29_2), .reg_weight21(reg_weight20_29_1), .reg_weight22(reg_weight20_29_2), .reg_activation12(reg_activation20_29_1), .reg_activation22(reg_activation20_29_2), .weight_en(weight_en));
SA22 U20_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_30_1), .partial_sum_in12(reg_psum19_30_2), .weight_in11(reg_weight19_30_1), .weight_in12(reg_weight19_30_2), .activation_in11(reg_activation20_29_1), .activation_in21(reg_activation20_29_2), .reg_partial_sum21(reg_psum20_30_1), .reg_partial_sum22(reg_psum20_30_2), .reg_weight21(reg_weight20_30_1), .reg_weight22(reg_weight20_30_2), .reg_activation12(reg_activation20_30_1), .reg_activation22(reg_activation20_30_2), .weight_en(weight_en));
SA22 U20_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_31_1), .partial_sum_in12(reg_psum19_31_2), .weight_in11(reg_weight19_31_1), .weight_in12(reg_weight19_31_2), .activation_in11(reg_activation20_30_1), .activation_in21(reg_activation20_30_2), .reg_partial_sum21(reg_psum20_31_1), .reg_partial_sum22(reg_psum20_31_2), .reg_weight21(reg_weight20_31_1), .reg_weight22(reg_weight20_31_2), .reg_activation12(reg_activation20_31_1), .reg_activation22(reg_activation20_31_2), .weight_en(weight_en));
SA22 U20_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum19_32_1), .partial_sum_in12(reg_psum19_32_2), .weight_in11(reg_weight19_32_1), .weight_in12(reg_weight19_32_2), .activation_in11(reg_activation20_31_1), .activation_in21(reg_activation20_31_2), .reg_partial_sum21(reg_psum20_32_1), .reg_partial_sum22(reg_psum20_32_2), .reg_weight21(reg_weight20_32_1), .reg_weight22(reg_weight20_32_2), .weight_en(weight_en));
SA22 U21_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_1_1), .partial_sum_in12(reg_psum20_1_2), .weight_in11(reg_weight20_1_1), .weight_in12(reg_weight20_1_2), .activation_in11(in_activation21_1_1), .activation_in21(in_activation21_1_2), .reg_partial_sum21(reg_psum21_1_1), .reg_partial_sum22(reg_psum21_1_2), .reg_weight21(reg_weight21_1_1), .reg_weight22(reg_weight21_1_2), .reg_activation12(reg_activation21_1_1), .reg_activation22(reg_activation21_1_2), .weight_en(weight_en));
SA22 U21_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_2_1), .partial_sum_in12(reg_psum20_2_2), .weight_in11(reg_weight20_2_1), .weight_in12(reg_weight20_2_2), .activation_in11(reg_activation21_1_1), .activation_in21(reg_activation21_1_2), .reg_partial_sum21(reg_psum21_2_1), .reg_partial_sum22(reg_psum21_2_2), .reg_weight21(reg_weight21_2_1), .reg_weight22(reg_weight21_2_2), .reg_activation12(reg_activation21_2_1), .reg_activation22(reg_activation21_2_2), .weight_en(weight_en));
SA22 U21_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_3_1), .partial_sum_in12(reg_psum20_3_2), .weight_in11(reg_weight20_3_1), .weight_in12(reg_weight20_3_2), .activation_in11(reg_activation21_2_1), .activation_in21(reg_activation21_2_2), .reg_partial_sum21(reg_psum21_3_1), .reg_partial_sum22(reg_psum21_3_2), .reg_weight21(reg_weight21_3_1), .reg_weight22(reg_weight21_3_2), .reg_activation12(reg_activation21_3_1), .reg_activation22(reg_activation21_3_2), .weight_en(weight_en));
SA22 U21_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_4_1), .partial_sum_in12(reg_psum20_4_2), .weight_in11(reg_weight20_4_1), .weight_in12(reg_weight20_4_2), .activation_in11(reg_activation21_3_1), .activation_in21(reg_activation21_3_2), .reg_partial_sum21(reg_psum21_4_1), .reg_partial_sum22(reg_psum21_4_2), .reg_weight21(reg_weight21_4_1), .reg_weight22(reg_weight21_4_2), .reg_activation12(reg_activation21_4_1), .reg_activation22(reg_activation21_4_2), .weight_en(weight_en));
SA22 U21_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_5_1), .partial_sum_in12(reg_psum20_5_2), .weight_in11(reg_weight20_5_1), .weight_in12(reg_weight20_5_2), .activation_in11(reg_activation21_4_1), .activation_in21(reg_activation21_4_2), .reg_partial_sum21(reg_psum21_5_1), .reg_partial_sum22(reg_psum21_5_2), .reg_weight21(reg_weight21_5_1), .reg_weight22(reg_weight21_5_2), .reg_activation12(reg_activation21_5_1), .reg_activation22(reg_activation21_5_2), .weight_en(weight_en));
SA22 U21_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_6_1), .partial_sum_in12(reg_psum20_6_2), .weight_in11(reg_weight20_6_1), .weight_in12(reg_weight20_6_2), .activation_in11(reg_activation21_5_1), .activation_in21(reg_activation21_5_2), .reg_partial_sum21(reg_psum21_6_1), .reg_partial_sum22(reg_psum21_6_2), .reg_weight21(reg_weight21_6_1), .reg_weight22(reg_weight21_6_2), .reg_activation12(reg_activation21_6_1), .reg_activation22(reg_activation21_6_2), .weight_en(weight_en));
SA22 U21_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_7_1), .partial_sum_in12(reg_psum20_7_2), .weight_in11(reg_weight20_7_1), .weight_in12(reg_weight20_7_2), .activation_in11(reg_activation21_6_1), .activation_in21(reg_activation21_6_2), .reg_partial_sum21(reg_psum21_7_1), .reg_partial_sum22(reg_psum21_7_2), .reg_weight21(reg_weight21_7_1), .reg_weight22(reg_weight21_7_2), .reg_activation12(reg_activation21_7_1), .reg_activation22(reg_activation21_7_2), .weight_en(weight_en));
SA22 U21_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_8_1), .partial_sum_in12(reg_psum20_8_2), .weight_in11(reg_weight20_8_1), .weight_in12(reg_weight20_8_2), .activation_in11(reg_activation21_7_1), .activation_in21(reg_activation21_7_2), .reg_partial_sum21(reg_psum21_8_1), .reg_partial_sum22(reg_psum21_8_2), .reg_weight21(reg_weight21_8_1), .reg_weight22(reg_weight21_8_2), .reg_activation12(reg_activation21_8_1), .reg_activation22(reg_activation21_8_2), .weight_en(weight_en));
SA22 U21_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_9_1), .partial_sum_in12(reg_psum20_9_2), .weight_in11(reg_weight20_9_1), .weight_in12(reg_weight20_9_2), .activation_in11(reg_activation21_8_1), .activation_in21(reg_activation21_8_2), .reg_partial_sum21(reg_psum21_9_1), .reg_partial_sum22(reg_psum21_9_2), .reg_weight21(reg_weight21_9_1), .reg_weight22(reg_weight21_9_2), .reg_activation12(reg_activation21_9_1), .reg_activation22(reg_activation21_9_2), .weight_en(weight_en));
SA22 U21_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_10_1), .partial_sum_in12(reg_psum20_10_2), .weight_in11(reg_weight20_10_1), .weight_in12(reg_weight20_10_2), .activation_in11(reg_activation21_9_1), .activation_in21(reg_activation21_9_2), .reg_partial_sum21(reg_psum21_10_1), .reg_partial_sum22(reg_psum21_10_2), .reg_weight21(reg_weight21_10_1), .reg_weight22(reg_weight21_10_2), .reg_activation12(reg_activation21_10_1), .reg_activation22(reg_activation21_10_2), .weight_en(weight_en));
SA22 U21_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_11_1), .partial_sum_in12(reg_psum20_11_2), .weight_in11(reg_weight20_11_1), .weight_in12(reg_weight20_11_2), .activation_in11(reg_activation21_10_1), .activation_in21(reg_activation21_10_2), .reg_partial_sum21(reg_psum21_11_1), .reg_partial_sum22(reg_psum21_11_2), .reg_weight21(reg_weight21_11_1), .reg_weight22(reg_weight21_11_2), .reg_activation12(reg_activation21_11_1), .reg_activation22(reg_activation21_11_2), .weight_en(weight_en));
SA22 U21_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_12_1), .partial_sum_in12(reg_psum20_12_2), .weight_in11(reg_weight20_12_1), .weight_in12(reg_weight20_12_2), .activation_in11(reg_activation21_11_1), .activation_in21(reg_activation21_11_2), .reg_partial_sum21(reg_psum21_12_1), .reg_partial_sum22(reg_psum21_12_2), .reg_weight21(reg_weight21_12_1), .reg_weight22(reg_weight21_12_2), .reg_activation12(reg_activation21_12_1), .reg_activation22(reg_activation21_12_2), .weight_en(weight_en));
SA22 U21_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_13_1), .partial_sum_in12(reg_psum20_13_2), .weight_in11(reg_weight20_13_1), .weight_in12(reg_weight20_13_2), .activation_in11(reg_activation21_12_1), .activation_in21(reg_activation21_12_2), .reg_partial_sum21(reg_psum21_13_1), .reg_partial_sum22(reg_psum21_13_2), .reg_weight21(reg_weight21_13_1), .reg_weight22(reg_weight21_13_2), .reg_activation12(reg_activation21_13_1), .reg_activation22(reg_activation21_13_2), .weight_en(weight_en));
SA22 U21_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_14_1), .partial_sum_in12(reg_psum20_14_2), .weight_in11(reg_weight20_14_1), .weight_in12(reg_weight20_14_2), .activation_in11(reg_activation21_13_1), .activation_in21(reg_activation21_13_2), .reg_partial_sum21(reg_psum21_14_1), .reg_partial_sum22(reg_psum21_14_2), .reg_weight21(reg_weight21_14_1), .reg_weight22(reg_weight21_14_2), .reg_activation12(reg_activation21_14_1), .reg_activation22(reg_activation21_14_2), .weight_en(weight_en));
SA22 U21_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_15_1), .partial_sum_in12(reg_psum20_15_2), .weight_in11(reg_weight20_15_1), .weight_in12(reg_weight20_15_2), .activation_in11(reg_activation21_14_1), .activation_in21(reg_activation21_14_2), .reg_partial_sum21(reg_psum21_15_1), .reg_partial_sum22(reg_psum21_15_2), .reg_weight21(reg_weight21_15_1), .reg_weight22(reg_weight21_15_2), .reg_activation12(reg_activation21_15_1), .reg_activation22(reg_activation21_15_2), .weight_en(weight_en));
SA22 U21_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_16_1), .partial_sum_in12(reg_psum20_16_2), .weight_in11(reg_weight20_16_1), .weight_in12(reg_weight20_16_2), .activation_in11(reg_activation21_15_1), .activation_in21(reg_activation21_15_2), .reg_partial_sum21(reg_psum21_16_1), .reg_partial_sum22(reg_psum21_16_2), .reg_weight21(reg_weight21_16_1), .reg_weight22(reg_weight21_16_2), .reg_activation12(reg_activation21_16_1), .reg_activation22(reg_activation21_16_2), .weight_en(weight_en));
SA22 U21_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_17_1), .partial_sum_in12(reg_psum20_17_2), .weight_in11(reg_weight20_17_1), .weight_in12(reg_weight20_17_2), .activation_in11(reg_activation21_16_1), .activation_in21(reg_activation21_16_2), .reg_partial_sum21(reg_psum21_17_1), .reg_partial_sum22(reg_psum21_17_2), .reg_weight21(reg_weight21_17_1), .reg_weight22(reg_weight21_17_2), .reg_activation12(reg_activation21_17_1), .reg_activation22(reg_activation21_17_2), .weight_en(weight_en));
SA22 U21_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_18_1), .partial_sum_in12(reg_psum20_18_2), .weight_in11(reg_weight20_18_1), .weight_in12(reg_weight20_18_2), .activation_in11(reg_activation21_17_1), .activation_in21(reg_activation21_17_2), .reg_partial_sum21(reg_psum21_18_1), .reg_partial_sum22(reg_psum21_18_2), .reg_weight21(reg_weight21_18_1), .reg_weight22(reg_weight21_18_2), .reg_activation12(reg_activation21_18_1), .reg_activation22(reg_activation21_18_2), .weight_en(weight_en));
SA22 U21_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_19_1), .partial_sum_in12(reg_psum20_19_2), .weight_in11(reg_weight20_19_1), .weight_in12(reg_weight20_19_2), .activation_in11(reg_activation21_18_1), .activation_in21(reg_activation21_18_2), .reg_partial_sum21(reg_psum21_19_1), .reg_partial_sum22(reg_psum21_19_2), .reg_weight21(reg_weight21_19_1), .reg_weight22(reg_weight21_19_2), .reg_activation12(reg_activation21_19_1), .reg_activation22(reg_activation21_19_2), .weight_en(weight_en));
SA22 U21_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_20_1), .partial_sum_in12(reg_psum20_20_2), .weight_in11(reg_weight20_20_1), .weight_in12(reg_weight20_20_2), .activation_in11(reg_activation21_19_1), .activation_in21(reg_activation21_19_2), .reg_partial_sum21(reg_psum21_20_1), .reg_partial_sum22(reg_psum21_20_2), .reg_weight21(reg_weight21_20_1), .reg_weight22(reg_weight21_20_2), .reg_activation12(reg_activation21_20_1), .reg_activation22(reg_activation21_20_2), .weight_en(weight_en));
SA22 U21_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_21_1), .partial_sum_in12(reg_psum20_21_2), .weight_in11(reg_weight20_21_1), .weight_in12(reg_weight20_21_2), .activation_in11(reg_activation21_20_1), .activation_in21(reg_activation21_20_2), .reg_partial_sum21(reg_psum21_21_1), .reg_partial_sum22(reg_psum21_21_2), .reg_weight21(reg_weight21_21_1), .reg_weight22(reg_weight21_21_2), .reg_activation12(reg_activation21_21_1), .reg_activation22(reg_activation21_21_2), .weight_en(weight_en));
SA22 U21_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_22_1), .partial_sum_in12(reg_psum20_22_2), .weight_in11(reg_weight20_22_1), .weight_in12(reg_weight20_22_2), .activation_in11(reg_activation21_21_1), .activation_in21(reg_activation21_21_2), .reg_partial_sum21(reg_psum21_22_1), .reg_partial_sum22(reg_psum21_22_2), .reg_weight21(reg_weight21_22_1), .reg_weight22(reg_weight21_22_2), .reg_activation12(reg_activation21_22_1), .reg_activation22(reg_activation21_22_2), .weight_en(weight_en));
SA22 U21_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_23_1), .partial_sum_in12(reg_psum20_23_2), .weight_in11(reg_weight20_23_1), .weight_in12(reg_weight20_23_2), .activation_in11(reg_activation21_22_1), .activation_in21(reg_activation21_22_2), .reg_partial_sum21(reg_psum21_23_1), .reg_partial_sum22(reg_psum21_23_2), .reg_weight21(reg_weight21_23_1), .reg_weight22(reg_weight21_23_2), .reg_activation12(reg_activation21_23_1), .reg_activation22(reg_activation21_23_2), .weight_en(weight_en));
SA22 U21_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_24_1), .partial_sum_in12(reg_psum20_24_2), .weight_in11(reg_weight20_24_1), .weight_in12(reg_weight20_24_2), .activation_in11(reg_activation21_23_1), .activation_in21(reg_activation21_23_2), .reg_partial_sum21(reg_psum21_24_1), .reg_partial_sum22(reg_psum21_24_2), .reg_weight21(reg_weight21_24_1), .reg_weight22(reg_weight21_24_2), .reg_activation12(reg_activation21_24_1), .reg_activation22(reg_activation21_24_2), .weight_en(weight_en));
SA22 U21_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_25_1), .partial_sum_in12(reg_psum20_25_2), .weight_in11(reg_weight20_25_1), .weight_in12(reg_weight20_25_2), .activation_in11(reg_activation21_24_1), .activation_in21(reg_activation21_24_2), .reg_partial_sum21(reg_psum21_25_1), .reg_partial_sum22(reg_psum21_25_2), .reg_weight21(reg_weight21_25_1), .reg_weight22(reg_weight21_25_2), .reg_activation12(reg_activation21_25_1), .reg_activation22(reg_activation21_25_2), .weight_en(weight_en));
SA22 U21_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_26_1), .partial_sum_in12(reg_psum20_26_2), .weight_in11(reg_weight20_26_1), .weight_in12(reg_weight20_26_2), .activation_in11(reg_activation21_25_1), .activation_in21(reg_activation21_25_2), .reg_partial_sum21(reg_psum21_26_1), .reg_partial_sum22(reg_psum21_26_2), .reg_weight21(reg_weight21_26_1), .reg_weight22(reg_weight21_26_2), .reg_activation12(reg_activation21_26_1), .reg_activation22(reg_activation21_26_2), .weight_en(weight_en));
SA22 U21_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_27_1), .partial_sum_in12(reg_psum20_27_2), .weight_in11(reg_weight20_27_1), .weight_in12(reg_weight20_27_2), .activation_in11(reg_activation21_26_1), .activation_in21(reg_activation21_26_2), .reg_partial_sum21(reg_psum21_27_1), .reg_partial_sum22(reg_psum21_27_2), .reg_weight21(reg_weight21_27_1), .reg_weight22(reg_weight21_27_2), .reg_activation12(reg_activation21_27_1), .reg_activation22(reg_activation21_27_2), .weight_en(weight_en));
SA22 U21_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_28_1), .partial_sum_in12(reg_psum20_28_2), .weight_in11(reg_weight20_28_1), .weight_in12(reg_weight20_28_2), .activation_in11(reg_activation21_27_1), .activation_in21(reg_activation21_27_2), .reg_partial_sum21(reg_psum21_28_1), .reg_partial_sum22(reg_psum21_28_2), .reg_weight21(reg_weight21_28_1), .reg_weight22(reg_weight21_28_2), .reg_activation12(reg_activation21_28_1), .reg_activation22(reg_activation21_28_2), .weight_en(weight_en));
SA22 U21_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_29_1), .partial_sum_in12(reg_psum20_29_2), .weight_in11(reg_weight20_29_1), .weight_in12(reg_weight20_29_2), .activation_in11(reg_activation21_28_1), .activation_in21(reg_activation21_28_2), .reg_partial_sum21(reg_psum21_29_1), .reg_partial_sum22(reg_psum21_29_2), .reg_weight21(reg_weight21_29_1), .reg_weight22(reg_weight21_29_2), .reg_activation12(reg_activation21_29_1), .reg_activation22(reg_activation21_29_2), .weight_en(weight_en));
SA22 U21_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_30_1), .partial_sum_in12(reg_psum20_30_2), .weight_in11(reg_weight20_30_1), .weight_in12(reg_weight20_30_2), .activation_in11(reg_activation21_29_1), .activation_in21(reg_activation21_29_2), .reg_partial_sum21(reg_psum21_30_1), .reg_partial_sum22(reg_psum21_30_2), .reg_weight21(reg_weight21_30_1), .reg_weight22(reg_weight21_30_2), .reg_activation12(reg_activation21_30_1), .reg_activation22(reg_activation21_30_2), .weight_en(weight_en));
SA22 U21_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_31_1), .partial_sum_in12(reg_psum20_31_2), .weight_in11(reg_weight20_31_1), .weight_in12(reg_weight20_31_2), .activation_in11(reg_activation21_30_1), .activation_in21(reg_activation21_30_2), .reg_partial_sum21(reg_psum21_31_1), .reg_partial_sum22(reg_psum21_31_2), .reg_weight21(reg_weight21_31_1), .reg_weight22(reg_weight21_31_2), .reg_activation12(reg_activation21_31_1), .reg_activation22(reg_activation21_31_2), .weight_en(weight_en));
SA22 U21_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum20_32_1), .partial_sum_in12(reg_psum20_32_2), .weight_in11(reg_weight20_32_1), .weight_in12(reg_weight20_32_2), .activation_in11(reg_activation21_31_1), .activation_in21(reg_activation21_31_2), .reg_partial_sum21(reg_psum21_32_1), .reg_partial_sum22(reg_psum21_32_2), .reg_weight21(reg_weight21_32_1), .reg_weight22(reg_weight21_32_2), .weight_en(weight_en));
SA22 U22_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_1_1), .partial_sum_in12(reg_psum21_1_2), .weight_in11(reg_weight21_1_1), .weight_in12(reg_weight21_1_2), .activation_in11(in_activation22_1_1), .activation_in21(in_activation22_1_2), .reg_partial_sum21(reg_psum22_1_1), .reg_partial_sum22(reg_psum22_1_2), .reg_weight21(reg_weight22_1_1), .reg_weight22(reg_weight22_1_2), .reg_activation12(reg_activation22_1_1), .reg_activation22(reg_activation22_1_2), .weight_en(weight_en));
SA22 U22_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_2_1), .partial_sum_in12(reg_psum21_2_2), .weight_in11(reg_weight21_2_1), .weight_in12(reg_weight21_2_2), .activation_in11(reg_activation22_1_1), .activation_in21(reg_activation22_1_2), .reg_partial_sum21(reg_psum22_2_1), .reg_partial_sum22(reg_psum22_2_2), .reg_weight21(reg_weight22_2_1), .reg_weight22(reg_weight22_2_2), .reg_activation12(reg_activation22_2_1), .reg_activation22(reg_activation22_2_2), .weight_en(weight_en));
SA22 U22_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_3_1), .partial_sum_in12(reg_psum21_3_2), .weight_in11(reg_weight21_3_1), .weight_in12(reg_weight21_3_2), .activation_in11(reg_activation22_2_1), .activation_in21(reg_activation22_2_2), .reg_partial_sum21(reg_psum22_3_1), .reg_partial_sum22(reg_psum22_3_2), .reg_weight21(reg_weight22_3_1), .reg_weight22(reg_weight22_3_2), .reg_activation12(reg_activation22_3_1), .reg_activation22(reg_activation22_3_2), .weight_en(weight_en));
SA22 U22_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_4_1), .partial_sum_in12(reg_psum21_4_2), .weight_in11(reg_weight21_4_1), .weight_in12(reg_weight21_4_2), .activation_in11(reg_activation22_3_1), .activation_in21(reg_activation22_3_2), .reg_partial_sum21(reg_psum22_4_1), .reg_partial_sum22(reg_psum22_4_2), .reg_weight21(reg_weight22_4_1), .reg_weight22(reg_weight22_4_2), .reg_activation12(reg_activation22_4_1), .reg_activation22(reg_activation22_4_2), .weight_en(weight_en));
SA22 U22_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_5_1), .partial_sum_in12(reg_psum21_5_2), .weight_in11(reg_weight21_5_1), .weight_in12(reg_weight21_5_2), .activation_in11(reg_activation22_4_1), .activation_in21(reg_activation22_4_2), .reg_partial_sum21(reg_psum22_5_1), .reg_partial_sum22(reg_psum22_5_2), .reg_weight21(reg_weight22_5_1), .reg_weight22(reg_weight22_5_2), .reg_activation12(reg_activation22_5_1), .reg_activation22(reg_activation22_5_2), .weight_en(weight_en));
SA22 U22_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_6_1), .partial_sum_in12(reg_psum21_6_2), .weight_in11(reg_weight21_6_1), .weight_in12(reg_weight21_6_2), .activation_in11(reg_activation22_5_1), .activation_in21(reg_activation22_5_2), .reg_partial_sum21(reg_psum22_6_1), .reg_partial_sum22(reg_psum22_6_2), .reg_weight21(reg_weight22_6_1), .reg_weight22(reg_weight22_6_2), .reg_activation12(reg_activation22_6_1), .reg_activation22(reg_activation22_6_2), .weight_en(weight_en));
SA22 U22_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_7_1), .partial_sum_in12(reg_psum21_7_2), .weight_in11(reg_weight21_7_1), .weight_in12(reg_weight21_7_2), .activation_in11(reg_activation22_6_1), .activation_in21(reg_activation22_6_2), .reg_partial_sum21(reg_psum22_7_1), .reg_partial_sum22(reg_psum22_7_2), .reg_weight21(reg_weight22_7_1), .reg_weight22(reg_weight22_7_2), .reg_activation12(reg_activation22_7_1), .reg_activation22(reg_activation22_7_2), .weight_en(weight_en));
SA22 U22_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_8_1), .partial_sum_in12(reg_psum21_8_2), .weight_in11(reg_weight21_8_1), .weight_in12(reg_weight21_8_2), .activation_in11(reg_activation22_7_1), .activation_in21(reg_activation22_7_2), .reg_partial_sum21(reg_psum22_8_1), .reg_partial_sum22(reg_psum22_8_2), .reg_weight21(reg_weight22_8_1), .reg_weight22(reg_weight22_8_2), .reg_activation12(reg_activation22_8_1), .reg_activation22(reg_activation22_8_2), .weight_en(weight_en));
SA22 U22_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_9_1), .partial_sum_in12(reg_psum21_9_2), .weight_in11(reg_weight21_9_1), .weight_in12(reg_weight21_9_2), .activation_in11(reg_activation22_8_1), .activation_in21(reg_activation22_8_2), .reg_partial_sum21(reg_psum22_9_1), .reg_partial_sum22(reg_psum22_9_2), .reg_weight21(reg_weight22_9_1), .reg_weight22(reg_weight22_9_2), .reg_activation12(reg_activation22_9_1), .reg_activation22(reg_activation22_9_2), .weight_en(weight_en));
SA22 U22_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_10_1), .partial_sum_in12(reg_psum21_10_2), .weight_in11(reg_weight21_10_1), .weight_in12(reg_weight21_10_2), .activation_in11(reg_activation22_9_1), .activation_in21(reg_activation22_9_2), .reg_partial_sum21(reg_psum22_10_1), .reg_partial_sum22(reg_psum22_10_2), .reg_weight21(reg_weight22_10_1), .reg_weight22(reg_weight22_10_2), .reg_activation12(reg_activation22_10_1), .reg_activation22(reg_activation22_10_2), .weight_en(weight_en));
SA22 U22_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_11_1), .partial_sum_in12(reg_psum21_11_2), .weight_in11(reg_weight21_11_1), .weight_in12(reg_weight21_11_2), .activation_in11(reg_activation22_10_1), .activation_in21(reg_activation22_10_2), .reg_partial_sum21(reg_psum22_11_1), .reg_partial_sum22(reg_psum22_11_2), .reg_weight21(reg_weight22_11_1), .reg_weight22(reg_weight22_11_2), .reg_activation12(reg_activation22_11_1), .reg_activation22(reg_activation22_11_2), .weight_en(weight_en));
SA22 U22_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_12_1), .partial_sum_in12(reg_psum21_12_2), .weight_in11(reg_weight21_12_1), .weight_in12(reg_weight21_12_2), .activation_in11(reg_activation22_11_1), .activation_in21(reg_activation22_11_2), .reg_partial_sum21(reg_psum22_12_1), .reg_partial_sum22(reg_psum22_12_2), .reg_weight21(reg_weight22_12_1), .reg_weight22(reg_weight22_12_2), .reg_activation12(reg_activation22_12_1), .reg_activation22(reg_activation22_12_2), .weight_en(weight_en));
SA22 U22_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_13_1), .partial_sum_in12(reg_psum21_13_2), .weight_in11(reg_weight21_13_1), .weight_in12(reg_weight21_13_2), .activation_in11(reg_activation22_12_1), .activation_in21(reg_activation22_12_2), .reg_partial_sum21(reg_psum22_13_1), .reg_partial_sum22(reg_psum22_13_2), .reg_weight21(reg_weight22_13_1), .reg_weight22(reg_weight22_13_2), .reg_activation12(reg_activation22_13_1), .reg_activation22(reg_activation22_13_2), .weight_en(weight_en));
SA22 U22_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_14_1), .partial_sum_in12(reg_psum21_14_2), .weight_in11(reg_weight21_14_1), .weight_in12(reg_weight21_14_2), .activation_in11(reg_activation22_13_1), .activation_in21(reg_activation22_13_2), .reg_partial_sum21(reg_psum22_14_1), .reg_partial_sum22(reg_psum22_14_2), .reg_weight21(reg_weight22_14_1), .reg_weight22(reg_weight22_14_2), .reg_activation12(reg_activation22_14_1), .reg_activation22(reg_activation22_14_2), .weight_en(weight_en));
SA22 U22_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_15_1), .partial_sum_in12(reg_psum21_15_2), .weight_in11(reg_weight21_15_1), .weight_in12(reg_weight21_15_2), .activation_in11(reg_activation22_14_1), .activation_in21(reg_activation22_14_2), .reg_partial_sum21(reg_psum22_15_1), .reg_partial_sum22(reg_psum22_15_2), .reg_weight21(reg_weight22_15_1), .reg_weight22(reg_weight22_15_2), .reg_activation12(reg_activation22_15_1), .reg_activation22(reg_activation22_15_2), .weight_en(weight_en));
SA22 U22_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_16_1), .partial_sum_in12(reg_psum21_16_2), .weight_in11(reg_weight21_16_1), .weight_in12(reg_weight21_16_2), .activation_in11(reg_activation22_15_1), .activation_in21(reg_activation22_15_2), .reg_partial_sum21(reg_psum22_16_1), .reg_partial_sum22(reg_psum22_16_2), .reg_weight21(reg_weight22_16_1), .reg_weight22(reg_weight22_16_2), .reg_activation12(reg_activation22_16_1), .reg_activation22(reg_activation22_16_2), .weight_en(weight_en));
SA22 U22_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_17_1), .partial_sum_in12(reg_psum21_17_2), .weight_in11(reg_weight21_17_1), .weight_in12(reg_weight21_17_2), .activation_in11(reg_activation22_16_1), .activation_in21(reg_activation22_16_2), .reg_partial_sum21(reg_psum22_17_1), .reg_partial_sum22(reg_psum22_17_2), .reg_weight21(reg_weight22_17_1), .reg_weight22(reg_weight22_17_2), .reg_activation12(reg_activation22_17_1), .reg_activation22(reg_activation22_17_2), .weight_en(weight_en));
SA22 U22_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_18_1), .partial_sum_in12(reg_psum21_18_2), .weight_in11(reg_weight21_18_1), .weight_in12(reg_weight21_18_2), .activation_in11(reg_activation22_17_1), .activation_in21(reg_activation22_17_2), .reg_partial_sum21(reg_psum22_18_1), .reg_partial_sum22(reg_psum22_18_2), .reg_weight21(reg_weight22_18_1), .reg_weight22(reg_weight22_18_2), .reg_activation12(reg_activation22_18_1), .reg_activation22(reg_activation22_18_2), .weight_en(weight_en));
SA22 U22_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_19_1), .partial_sum_in12(reg_psum21_19_2), .weight_in11(reg_weight21_19_1), .weight_in12(reg_weight21_19_2), .activation_in11(reg_activation22_18_1), .activation_in21(reg_activation22_18_2), .reg_partial_sum21(reg_psum22_19_1), .reg_partial_sum22(reg_psum22_19_2), .reg_weight21(reg_weight22_19_1), .reg_weight22(reg_weight22_19_2), .reg_activation12(reg_activation22_19_1), .reg_activation22(reg_activation22_19_2), .weight_en(weight_en));
SA22 U22_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_20_1), .partial_sum_in12(reg_psum21_20_2), .weight_in11(reg_weight21_20_1), .weight_in12(reg_weight21_20_2), .activation_in11(reg_activation22_19_1), .activation_in21(reg_activation22_19_2), .reg_partial_sum21(reg_psum22_20_1), .reg_partial_sum22(reg_psum22_20_2), .reg_weight21(reg_weight22_20_1), .reg_weight22(reg_weight22_20_2), .reg_activation12(reg_activation22_20_1), .reg_activation22(reg_activation22_20_2), .weight_en(weight_en));
SA22 U22_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_21_1), .partial_sum_in12(reg_psum21_21_2), .weight_in11(reg_weight21_21_1), .weight_in12(reg_weight21_21_2), .activation_in11(reg_activation22_20_1), .activation_in21(reg_activation22_20_2), .reg_partial_sum21(reg_psum22_21_1), .reg_partial_sum22(reg_psum22_21_2), .reg_weight21(reg_weight22_21_1), .reg_weight22(reg_weight22_21_2), .reg_activation12(reg_activation22_21_1), .reg_activation22(reg_activation22_21_2), .weight_en(weight_en));
SA22 U22_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_22_1), .partial_sum_in12(reg_psum21_22_2), .weight_in11(reg_weight21_22_1), .weight_in12(reg_weight21_22_2), .activation_in11(reg_activation22_21_1), .activation_in21(reg_activation22_21_2), .reg_partial_sum21(reg_psum22_22_1), .reg_partial_sum22(reg_psum22_22_2), .reg_weight21(reg_weight22_22_1), .reg_weight22(reg_weight22_22_2), .reg_activation12(reg_activation22_22_1), .reg_activation22(reg_activation22_22_2), .weight_en(weight_en));
SA22 U22_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_23_1), .partial_sum_in12(reg_psum21_23_2), .weight_in11(reg_weight21_23_1), .weight_in12(reg_weight21_23_2), .activation_in11(reg_activation22_22_1), .activation_in21(reg_activation22_22_2), .reg_partial_sum21(reg_psum22_23_1), .reg_partial_sum22(reg_psum22_23_2), .reg_weight21(reg_weight22_23_1), .reg_weight22(reg_weight22_23_2), .reg_activation12(reg_activation22_23_1), .reg_activation22(reg_activation22_23_2), .weight_en(weight_en));
SA22 U22_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_24_1), .partial_sum_in12(reg_psum21_24_2), .weight_in11(reg_weight21_24_1), .weight_in12(reg_weight21_24_2), .activation_in11(reg_activation22_23_1), .activation_in21(reg_activation22_23_2), .reg_partial_sum21(reg_psum22_24_1), .reg_partial_sum22(reg_psum22_24_2), .reg_weight21(reg_weight22_24_1), .reg_weight22(reg_weight22_24_2), .reg_activation12(reg_activation22_24_1), .reg_activation22(reg_activation22_24_2), .weight_en(weight_en));
SA22 U22_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_25_1), .partial_sum_in12(reg_psum21_25_2), .weight_in11(reg_weight21_25_1), .weight_in12(reg_weight21_25_2), .activation_in11(reg_activation22_24_1), .activation_in21(reg_activation22_24_2), .reg_partial_sum21(reg_psum22_25_1), .reg_partial_sum22(reg_psum22_25_2), .reg_weight21(reg_weight22_25_1), .reg_weight22(reg_weight22_25_2), .reg_activation12(reg_activation22_25_1), .reg_activation22(reg_activation22_25_2), .weight_en(weight_en));
SA22 U22_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_26_1), .partial_sum_in12(reg_psum21_26_2), .weight_in11(reg_weight21_26_1), .weight_in12(reg_weight21_26_2), .activation_in11(reg_activation22_25_1), .activation_in21(reg_activation22_25_2), .reg_partial_sum21(reg_psum22_26_1), .reg_partial_sum22(reg_psum22_26_2), .reg_weight21(reg_weight22_26_1), .reg_weight22(reg_weight22_26_2), .reg_activation12(reg_activation22_26_1), .reg_activation22(reg_activation22_26_2), .weight_en(weight_en));
SA22 U22_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_27_1), .partial_sum_in12(reg_psum21_27_2), .weight_in11(reg_weight21_27_1), .weight_in12(reg_weight21_27_2), .activation_in11(reg_activation22_26_1), .activation_in21(reg_activation22_26_2), .reg_partial_sum21(reg_psum22_27_1), .reg_partial_sum22(reg_psum22_27_2), .reg_weight21(reg_weight22_27_1), .reg_weight22(reg_weight22_27_2), .reg_activation12(reg_activation22_27_1), .reg_activation22(reg_activation22_27_2), .weight_en(weight_en));
SA22 U22_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_28_1), .partial_sum_in12(reg_psum21_28_2), .weight_in11(reg_weight21_28_1), .weight_in12(reg_weight21_28_2), .activation_in11(reg_activation22_27_1), .activation_in21(reg_activation22_27_2), .reg_partial_sum21(reg_psum22_28_1), .reg_partial_sum22(reg_psum22_28_2), .reg_weight21(reg_weight22_28_1), .reg_weight22(reg_weight22_28_2), .reg_activation12(reg_activation22_28_1), .reg_activation22(reg_activation22_28_2), .weight_en(weight_en));
SA22 U22_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_29_1), .partial_sum_in12(reg_psum21_29_2), .weight_in11(reg_weight21_29_1), .weight_in12(reg_weight21_29_2), .activation_in11(reg_activation22_28_1), .activation_in21(reg_activation22_28_2), .reg_partial_sum21(reg_psum22_29_1), .reg_partial_sum22(reg_psum22_29_2), .reg_weight21(reg_weight22_29_1), .reg_weight22(reg_weight22_29_2), .reg_activation12(reg_activation22_29_1), .reg_activation22(reg_activation22_29_2), .weight_en(weight_en));
SA22 U22_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_30_1), .partial_sum_in12(reg_psum21_30_2), .weight_in11(reg_weight21_30_1), .weight_in12(reg_weight21_30_2), .activation_in11(reg_activation22_29_1), .activation_in21(reg_activation22_29_2), .reg_partial_sum21(reg_psum22_30_1), .reg_partial_sum22(reg_psum22_30_2), .reg_weight21(reg_weight22_30_1), .reg_weight22(reg_weight22_30_2), .reg_activation12(reg_activation22_30_1), .reg_activation22(reg_activation22_30_2), .weight_en(weight_en));
SA22 U22_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_31_1), .partial_sum_in12(reg_psum21_31_2), .weight_in11(reg_weight21_31_1), .weight_in12(reg_weight21_31_2), .activation_in11(reg_activation22_30_1), .activation_in21(reg_activation22_30_2), .reg_partial_sum21(reg_psum22_31_1), .reg_partial_sum22(reg_psum22_31_2), .reg_weight21(reg_weight22_31_1), .reg_weight22(reg_weight22_31_2), .reg_activation12(reg_activation22_31_1), .reg_activation22(reg_activation22_31_2), .weight_en(weight_en));
SA22 U22_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum21_32_1), .partial_sum_in12(reg_psum21_32_2), .weight_in11(reg_weight21_32_1), .weight_in12(reg_weight21_32_2), .activation_in11(reg_activation22_31_1), .activation_in21(reg_activation22_31_2), .reg_partial_sum21(reg_psum22_32_1), .reg_partial_sum22(reg_psum22_32_2), .reg_weight21(reg_weight22_32_1), .reg_weight22(reg_weight22_32_2), .weight_en(weight_en));
SA22 U23_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_1_1), .partial_sum_in12(reg_psum22_1_2), .weight_in11(reg_weight22_1_1), .weight_in12(reg_weight22_1_2), .activation_in11(in_activation23_1_1), .activation_in21(in_activation23_1_2), .reg_partial_sum21(reg_psum23_1_1), .reg_partial_sum22(reg_psum23_1_2), .reg_weight21(reg_weight23_1_1), .reg_weight22(reg_weight23_1_2), .reg_activation12(reg_activation23_1_1), .reg_activation22(reg_activation23_1_2), .weight_en(weight_en));
SA22 U23_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_2_1), .partial_sum_in12(reg_psum22_2_2), .weight_in11(reg_weight22_2_1), .weight_in12(reg_weight22_2_2), .activation_in11(reg_activation23_1_1), .activation_in21(reg_activation23_1_2), .reg_partial_sum21(reg_psum23_2_1), .reg_partial_sum22(reg_psum23_2_2), .reg_weight21(reg_weight23_2_1), .reg_weight22(reg_weight23_2_2), .reg_activation12(reg_activation23_2_1), .reg_activation22(reg_activation23_2_2), .weight_en(weight_en));
SA22 U23_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_3_1), .partial_sum_in12(reg_psum22_3_2), .weight_in11(reg_weight22_3_1), .weight_in12(reg_weight22_3_2), .activation_in11(reg_activation23_2_1), .activation_in21(reg_activation23_2_2), .reg_partial_sum21(reg_psum23_3_1), .reg_partial_sum22(reg_psum23_3_2), .reg_weight21(reg_weight23_3_1), .reg_weight22(reg_weight23_3_2), .reg_activation12(reg_activation23_3_1), .reg_activation22(reg_activation23_3_2), .weight_en(weight_en));
SA22 U23_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_4_1), .partial_sum_in12(reg_psum22_4_2), .weight_in11(reg_weight22_4_1), .weight_in12(reg_weight22_4_2), .activation_in11(reg_activation23_3_1), .activation_in21(reg_activation23_3_2), .reg_partial_sum21(reg_psum23_4_1), .reg_partial_sum22(reg_psum23_4_2), .reg_weight21(reg_weight23_4_1), .reg_weight22(reg_weight23_4_2), .reg_activation12(reg_activation23_4_1), .reg_activation22(reg_activation23_4_2), .weight_en(weight_en));
SA22 U23_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_5_1), .partial_sum_in12(reg_psum22_5_2), .weight_in11(reg_weight22_5_1), .weight_in12(reg_weight22_5_2), .activation_in11(reg_activation23_4_1), .activation_in21(reg_activation23_4_2), .reg_partial_sum21(reg_psum23_5_1), .reg_partial_sum22(reg_psum23_5_2), .reg_weight21(reg_weight23_5_1), .reg_weight22(reg_weight23_5_2), .reg_activation12(reg_activation23_5_1), .reg_activation22(reg_activation23_5_2), .weight_en(weight_en));
SA22 U23_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_6_1), .partial_sum_in12(reg_psum22_6_2), .weight_in11(reg_weight22_6_1), .weight_in12(reg_weight22_6_2), .activation_in11(reg_activation23_5_1), .activation_in21(reg_activation23_5_2), .reg_partial_sum21(reg_psum23_6_1), .reg_partial_sum22(reg_psum23_6_2), .reg_weight21(reg_weight23_6_1), .reg_weight22(reg_weight23_6_2), .reg_activation12(reg_activation23_6_1), .reg_activation22(reg_activation23_6_2), .weight_en(weight_en));
SA22 U23_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_7_1), .partial_sum_in12(reg_psum22_7_2), .weight_in11(reg_weight22_7_1), .weight_in12(reg_weight22_7_2), .activation_in11(reg_activation23_6_1), .activation_in21(reg_activation23_6_2), .reg_partial_sum21(reg_psum23_7_1), .reg_partial_sum22(reg_psum23_7_2), .reg_weight21(reg_weight23_7_1), .reg_weight22(reg_weight23_7_2), .reg_activation12(reg_activation23_7_1), .reg_activation22(reg_activation23_7_2), .weight_en(weight_en));
SA22 U23_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_8_1), .partial_sum_in12(reg_psum22_8_2), .weight_in11(reg_weight22_8_1), .weight_in12(reg_weight22_8_2), .activation_in11(reg_activation23_7_1), .activation_in21(reg_activation23_7_2), .reg_partial_sum21(reg_psum23_8_1), .reg_partial_sum22(reg_psum23_8_2), .reg_weight21(reg_weight23_8_1), .reg_weight22(reg_weight23_8_2), .reg_activation12(reg_activation23_8_1), .reg_activation22(reg_activation23_8_2), .weight_en(weight_en));
SA22 U23_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_9_1), .partial_sum_in12(reg_psum22_9_2), .weight_in11(reg_weight22_9_1), .weight_in12(reg_weight22_9_2), .activation_in11(reg_activation23_8_1), .activation_in21(reg_activation23_8_2), .reg_partial_sum21(reg_psum23_9_1), .reg_partial_sum22(reg_psum23_9_2), .reg_weight21(reg_weight23_9_1), .reg_weight22(reg_weight23_9_2), .reg_activation12(reg_activation23_9_1), .reg_activation22(reg_activation23_9_2), .weight_en(weight_en));
SA22 U23_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_10_1), .partial_sum_in12(reg_psum22_10_2), .weight_in11(reg_weight22_10_1), .weight_in12(reg_weight22_10_2), .activation_in11(reg_activation23_9_1), .activation_in21(reg_activation23_9_2), .reg_partial_sum21(reg_psum23_10_1), .reg_partial_sum22(reg_psum23_10_2), .reg_weight21(reg_weight23_10_1), .reg_weight22(reg_weight23_10_2), .reg_activation12(reg_activation23_10_1), .reg_activation22(reg_activation23_10_2), .weight_en(weight_en));
SA22 U23_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_11_1), .partial_sum_in12(reg_psum22_11_2), .weight_in11(reg_weight22_11_1), .weight_in12(reg_weight22_11_2), .activation_in11(reg_activation23_10_1), .activation_in21(reg_activation23_10_2), .reg_partial_sum21(reg_psum23_11_1), .reg_partial_sum22(reg_psum23_11_2), .reg_weight21(reg_weight23_11_1), .reg_weight22(reg_weight23_11_2), .reg_activation12(reg_activation23_11_1), .reg_activation22(reg_activation23_11_2), .weight_en(weight_en));
SA22 U23_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_12_1), .partial_sum_in12(reg_psum22_12_2), .weight_in11(reg_weight22_12_1), .weight_in12(reg_weight22_12_2), .activation_in11(reg_activation23_11_1), .activation_in21(reg_activation23_11_2), .reg_partial_sum21(reg_psum23_12_1), .reg_partial_sum22(reg_psum23_12_2), .reg_weight21(reg_weight23_12_1), .reg_weight22(reg_weight23_12_2), .reg_activation12(reg_activation23_12_1), .reg_activation22(reg_activation23_12_2), .weight_en(weight_en));
SA22 U23_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_13_1), .partial_sum_in12(reg_psum22_13_2), .weight_in11(reg_weight22_13_1), .weight_in12(reg_weight22_13_2), .activation_in11(reg_activation23_12_1), .activation_in21(reg_activation23_12_2), .reg_partial_sum21(reg_psum23_13_1), .reg_partial_sum22(reg_psum23_13_2), .reg_weight21(reg_weight23_13_1), .reg_weight22(reg_weight23_13_2), .reg_activation12(reg_activation23_13_1), .reg_activation22(reg_activation23_13_2), .weight_en(weight_en));
SA22 U23_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_14_1), .partial_sum_in12(reg_psum22_14_2), .weight_in11(reg_weight22_14_1), .weight_in12(reg_weight22_14_2), .activation_in11(reg_activation23_13_1), .activation_in21(reg_activation23_13_2), .reg_partial_sum21(reg_psum23_14_1), .reg_partial_sum22(reg_psum23_14_2), .reg_weight21(reg_weight23_14_1), .reg_weight22(reg_weight23_14_2), .reg_activation12(reg_activation23_14_1), .reg_activation22(reg_activation23_14_2), .weight_en(weight_en));
SA22 U23_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_15_1), .partial_sum_in12(reg_psum22_15_2), .weight_in11(reg_weight22_15_1), .weight_in12(reg_weight22_15_2), .activation_in11(reg_activation23_14_1), .activation_in21(reg_activation23_14_2), .reg_partial_sum21(reg_psum23_15_1), .reg_partial_sum22(reg_psum23_15_2), .reg_weight21(reg_weight23_15_1), .reg_weight22(reg_weight23_15_2), .reg_activation12(reg_activation23_15_1), .reg_activation22(reg_activation23_15_2), .weight_en(weight_en));
SA22 U23_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_16_1), .partial_sum_in12(reg_psum22_16_2), .weight_in11(reg_weight22_16_1), .weight_in12(reg_weight22_16_2), .activation_in11(reg_activation23_15_1), .activation_in21(reg_activation23_15_2), .reg_partial_sum21(reg_psum23_16_1), .reg_partial_sum22(reg_psum23_16_2), .reg_weight21(reg_weight23_16_1), .reg_weight22(reg_weight23_16_2), .reg_activation12(reg_activation23_16_1), .reg_activation22(reg_activation23_16_2), .weight_en(weight_en));
SA22 U23_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_17_1), .partial_sum_in12(reg_psum22_17_2), .weight_in11(reg_weight22_17_1), .weight_in12(reg_weight22_17_2), .activation_in11(reg_activation23_16_1), .activation_in21(reg_activation23_16_2), .reg_partial_sum21(reg_psum23_17_1), .reg_partial_sum22(reg_psum23_17_2), .reg_weight21(reg_weight23_17_1), .reg_weight22(reg_weight23_17_2), .reg_activation12(reg_activation23_17_1), .reg_activation22(reg_activation23_17_2), .weight_en(weight_en));
SA22 U23_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_18_1), .partial_sum_in12(reg_psum22_18_2), .weight_in11(reg_weight22_18_1), .weight_in12(reg_weight22_18_2), .activation_in11(reg_activation23_17_1), .activation_in21(reg_activation23_17_2), .reg_partial_sum21(reg_psum23_18_1), .reg_partial_sum22(reg_psum23_18_2), .reg_weight21(reg_weight23_18_1), .reg_weight22(reg_weight23_18_2), .reg_activation12(reg_activation23_18_1), .reg_activation22(reg_activation23_18_2), .weight_en(weight_en));
SA22 U23_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_19_1), .partial_sum_in12(reg_psum22_19_2), .weight_in11(reg_weight22_19_1), .weight_in12(reg_weight22_19_2), .activation_in11(reg_activation23_18_1), .activation_in21(reg_activation23_18_2), .reg_partial_sum21(reg_psum23_19_1), .reg_partial_sum22(reg_psum23_19_2), .reg_weight21(reg_weight23_19_1), .reg_weight22(reg_weight23_19_2), .reg_activation12(reg_activation23_19_1), .reg_activation22(reg_activation23_19_2), .weight_en(weight_en));
SA22 U23_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_20_1), .partial_sum_in12(reg_psum22_20_2), .weight_in11(reg_weight22_20_1), .weight_in12(reg_weight22_20_2), .activation_in11(reg_activation23_19_1), .activation_in21(reg_activation23_19_2), .reg_partial_sum21(reg_psum23_20_1), .reg_partial_sum22(reg_psum23_20_2), .reg_weight21(reg_weight23_20_1), .reg_weight22(reg_weight23_20_2), .reg_activation12(reg_activation23_20_1), .reg_activation22(reg_activation23_20_2), .weight_en(weight_en));
SA22 U23_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_21_1), .partial_sum_in12(reg_psum22_21_2), .weight_in11(reg_weight22_21_1), .weight_in12(reg_weight22_21_2), .activation_in11(reg_activation23_20_1), .activation_in21(reg_activation23_20_2), .reg_partial_sum21(reg_psum23_21_1), .reg_partial_sum22(reg_psum23_21_2), .reg_weight21(reg_weight23_21_1), .reg_weight22(reg_weight23_21_2), .reg_activation12(reg_activation23_21_1), .reg_activation22(reg_activation23_21_2), .weight_en(weight_en));
SA22 U23_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_22_1), .partial_sum_in12(reg_psum22_22_2), .weight_in11(reg_weight22_22_1), .weight_in12(reg_weight22_22_2), .activation_in11(reg_activation23_21_1), .activation_in21(reg_activation23_21_2), .reg_partial_sum21(reg_psum23_22_1), .reg_partial_sum22(reg_psum23_22_2), .reg_weight21(reg_weight23_22_1), .reg_weight22(reg_weight23_22_2), .reg_activation12(reg_activation23_22_1), .reg_activation22(reg_activation23_22_2), .weight_en(weight_en));
SA22 U23_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_23_1), .partial_sum_in12(reg_psum22_23_2), .weight_in11(reg_weight22_23_1), .weight_in12(reg_weight22_23_2), .activation_in11(reg_activation23_22_1), .activation_in21(reg_activation23_22_2), .reg_partial_sum21(reg_psum23_23_1), .reg_partial_sum22(reg_psum23_23_2), .reg_weight21(reg_weight23_23_1), .reg_weight22(reg_weight23_23_2), .reg_activation12(reg_activation23_23_1), .reg_activation22(reg_activation23_23_2), .weight_en(weight_en));
SA22 U23_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_24_1), .partial_sum_in12(reg_psum22_24_2), .weight_in11(reg_weight22_24_1), .weight_in12(reg_weight22_24_2), .activation_in11(reg_activation23_23_1), .activation_in21(reg_activation23_23_2), .reg_partial_sum21(reg_psum23_24_1), .reg_partial_sum22(reg_psum23_24_2), .reg_weight21(reg_weight23_24_1), .reg_weight22(reg_weight23_24_2), .reg_activation12(reg_activation23_24_1), .reg_activation22(reg_activation23_24_2), .weight_en(weight_en));
SA22 U23_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_25_1), .partial_sum_in12(reg_psum22_25_2), .weight_in11(reg_weight22_25_1), .weight_in12(reg_weight22_25_2), .activation_in11(reg_activation23_24_1), .activation_in21(reg_activation23_24_2), .reg_partial_sum21(reg_psum23_25_1), .reg_partial_sum22(reg_psum23_25_2), .reg_weight21(reg_weight23_25_1), .reg_weight22(reg_weight23_25_2), .reg_activation12(reg_activation23_25_1), .reg_activation22(reg_activation23_25_2), .weight_en(weight_en));
SA22 U23_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_26_1), .partial_sum_in12(reg_psum22_26_2), .weight_in11(reg_weight22_26_1), .weight_in12(reg_weight22_26_2), .activation_in11(reg_activation23_25_1), .activation_in21(reg_activation23_25_2), .reg_partial_sum21(reg_psum23_26_1), .reg_partial_sum22(reg_psum23_26_2), .reg_weight21(reg_weight23_26_1), .reg_weight22(reg_weight23_26_2), .reg_activation12(reg_activation23_26_1), .reg_activation22(reg_activation23_26_2), .weight_en(weight_en));
SA22 U23_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_27_1), .partial_sum_in12(reg_psum22_27_2), .weight_in11(reg_weight22_27_1), .weight_in12(reg_weight22_27_2), .activation_in11(reg_activation23_26_1), .activation_in21(reg_activation23_26_2), .reg_partial_sum21(reg_psum23_27_1), .reg_partial_sum22(reg_psum23_27_2), .reg_weight21(reg_weight23_27_1), .reg_weight22(reg_weight23_27_2), .reg_activation12(reg_activation23_27_1), .reg_activation22(reg_activation23_27_2), .weight_en(weight_en));
SA22 U23_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_28_1), .partial_sum_in12(reg_psum22_28_2), .weight_in11(reg_weight22_28_1), .weight_in12(reg_weight22_28_2), .activation_in11(reg_activation23_27_1), .activation_in21(reg_activation23_27_2), .reg_partial_sum21(reg_psum23_28_1), .reg_partial_sum22(reg_psum23_28_2), .reg_weight21(reg_weight23_28_1), .reg_weight22(reg_weight23_28_2), .reg_activation12(reg_activation23_28_1), .reg_activation22(reg_activation23_28_2), .weight_en(weight_en));
SA22 U23_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_29_1), .partial_sum_in12(reg_psum22_29_2), .weight_in11(reg_weight22_29_1), .weight_in12(reg_weight22_29_2), .activation_in11(reg_activation23_28_1), .activation_in21(reg_activation23_28_2), .reg_partial_sum21(reg_psum23_29_1), .reg_partial_sum22(reg_psum23_29_2), .reg_weight21(reg_weight23_29_1), .reg_weight22(reg_weight23_29_2), .reg_activation12(reg_activation23_29_1), .reg_activation22(reg_activation23_29_2), .weight_en(weight_en));
SA22 U23_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_30_1), .partial_sum_in12(reg_psum22_30_2), .weight_in11(reg_weight22_30_1), .weight_in12(reg_weight22_30_2), .activation_in11(reg_activation23_29_1), .activation_in21(reg_activation23_29_2), .reg_partial_sum21(reg_psum23_30_1), .reg_partial_sum22(reg_psum23_30_2), .reg_weight21(reg_weight23_30_1), .reg_weight22(reg_weight23_30_2), .reg_activation12(reg_activation23_30_1), .reg_activation22(reg_activation23_30_2), .weight_en(weight_en));
SA22 U23_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_31_1), .partial_sum_in12(reg_psum22_31_2), .weight_in11(reg_weight22_31_1), .weight_in12(reg_weight22_31_2), .activation_in11(reg_activation23_30_1), .activation_in21(reg_activation23_30_2), .reg_partial_sum21(reg_psum23_31_1), .reg_partial_sum22(reg_psum23_31_2), .reg_weight21(reg_weight23_31_1), .reg_weight22(reg_weight23_31_2), .reg_activation12(reg_activation23_31_1), .reg_activation22(reg_activation23_31_2), .weight_en(weight_en));
SA22 U23_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum22_32_1), .partial_sum_in12(reg_psum22_32_2), .weight_in11(reg_weight22_32_1), .weight_in12(reg_weight22_32_2), .activation_in11(reg_activation23_31_1), .activation_in21(reg_activation23_31_2), .reg_partial_sum21(reg_psum23_32_1), .reg_partial_sum22(reg_psum23_32_2), .reg_weight21(reg_weight23_32_1), .reg_weight22(reg_weight23_32_2), .weight_en(weight_en));
SA22 U24_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_1_1), .partial_sum_in12(reg_psum23_1_2), .weight_in11(reg_weight23_1_1), .weight_in12(reg_weight23_1_2), .activation_in11(in_activation24_1_1), .activation_in21(in_activation24_1_2), .reg_partial_sum21(reg_psum24_1_1), .reg_partial_sum22(reg_psum24_1_2), .reg_weight21(reg_weight24_1_1), .reg_weight22(reg_weight24_1_2), .reg_activation12(reg_activation24_1_1), .reg_activation22(reg_activation24_1_2), .weight_en(weight_en));
SA22 U24_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_2_1), .partial_sum_in12(reg_psum23_2_2), .weight_in11(reg_weight23_2_1), .weight_in12(reg_weight23_2_2), .activation_in11(reg_activation24_1_1), .activation_in21(reg_activation24_1_2), .reg_partial_sum21(reg_psum24_2_1), .reg_partial_sum22(reg_psum24_2_2), .reg_weight21(reg_weight24_2_1), .reg_weight22(reg_weight24_2_2), .reg_activation12(reg_activation24_2_1), .reg_activation22(reg_activation24_2_2), .weight_en(weight_en));
SA22 U24_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_3_1), .partial_sum_in12(reg_psum23_3_2), .weight_in11(reg_weight23_3_1), .weight_in12(reg_weight23_3_2), .activation_in11(reg_activation24_2_1), .activation_in21(reg_activation24_2_2), .reg_partial_sum21(reg_psum24_3_1), .reg_partial_sum22(reg_psum24_3_2), .reg_weight21(reg_weight24_3_1), .reg_weight22(reg_weight24_3_2), .reg_activation12(reg_activation24_3_1), .reg_activation22(reg_activation24_3_2), .weight_en(weight_en));
SA22 U24_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_4_1), .partial_sum_in12(reg_psum23_4_2), .weight_in11(reg_weight23_4_1), .weight_in12(reg_weight23_4_2), .activation_in11(reg_activation24_3_1), .activation_in21(reg_activation24_3_2), .reg_partial_sum21(reg_psum24_4_1), .reg_partial_sum22(reg_psum24_4_2), .reg_weight21(reg_weight24_4_1), .reg_weight22(reg_weight24_4_2), .reg_activation12(reg_activation24_4_1), .reg_activation22(reg_activation24_4_2), .weight_en(weight_en));
SA22 U24_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_5_1), .partial_sum_in12(reg_psum23_5_2), .weight_in11(reg_weight23_5_1), .weight_in12(reg_weight23_5_2), .activation_in11(reg_activation24_4_1), .activation_in21(reg_activation24_4_2), .reg_partial_sum21(reg_psum24_5_1), .reg_partial_sum22(reg_psum24_5_2), .reg_weight21(reg_weight24_5_1), .reg_weight22(reg_weight24_5_2), .reg_activation12(reg_activation24_5_1), .reg_activation22(reg_activation24_5_2), .weight_en(weight_en));
SA22 U24_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_6_1), .partial_sum_in12(reg_psum23_6_2), .weight_in11(reg_weight23_6_1), .weight_in12(reg_weight23_6_2), .activation_in11(reg_activation24_5_1), .activation_in21(reg_activation24_5_2), .reg_partial_sum21(reg_psum24_6_1), .reg_partial_sum22(reg_psum24_6_2), .reg_weight21(reg_weight24_6_1), .reg_weight22(reg_weight24_6_2), .reg_activation12(reg_activation24_6_1), .reg_activation22(reg_activation24_6_2), .weight_en(weight_en));
SA22 U24_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_7_1), .partial_sum_in12(reg_psum23_7_2), .weight_in11(reg_weight23_7_1), .weight_in12(reg_weight23_7_2), .activation_in11(reg_activation24_6_1), .activation_in21(reg_activation24_6_2), .reg_partial_sum21(reg_psum24_7_1), .reg_partial_sum22(reg_psum24_7_2), .reg_weight21(reg_weight24_7_1), .reg_weight22(reg_weight24_7_2), .reg_activation12(reg_activation24_7_1), .reg_activation22(reg_activation24_7_2), .weight_en(weight_en));
SA22 U24_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_8_1), .partial_sum_in12(reg_psum23_8_2), .weight_in11(reg_weight23_8_1), .weight_in12(reg_weight23_8_2), .activation_in11(reg_activation24_7_1), .activation_in21(reg_activation24_7_2), .reg_partial_sum21(reg_psum24_8_1), .reg_partial_sum22(reg_psum24_8_2), .reg_weight21(reg_weight24_8_1), .reg_weight22(reg_weight24_8_2), .reg_activation12(reg_activation24_8_1), .reg_activation22(reg_activation24_8_2), .weight_en(weight_en));
SA22 U24_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_9_1), .partial_sum_in12(reg_psum23_9_2), .weight_in11(reg_weight23_9_1), .weight_in12(reg_weight23_9_2), .activation_in11(reg_activation24_8_1), .activation_in21(reg_activation24_8_2), .reg_partial_sum21(reg_psum24_9_1), .reg_partial_sum22(reg_psum24_9_2), .reg_weight21(reg_weight24_9_1), .reg_weight22(reg_weight24_9_2), .reg_activation12(reg_activation24_9_1), .reg_activation22(reg_activation24_9_2), .weight_en(weight_en));
SA22 U24_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_10_1), .partial_sum_in12(reg_psum23_10_2), .weight_in11(reg_weight23_10_1), .weight_in12(reg_weight23_10_2), .activation_in11(reg_activation24_9_1), .activation_in21(reg_activation24_9_2), .reg_partial_sum21(reg_psum24_10_1), .reg_partial_sum22(reg_psum24_10_2), .reg_weight21(reg_weight24_10_1), .reg_weight22(reg_weight24_10_2), .reg_activation12(reg_activation24_10_1), .reg_activation22(reg_activation24_10_2), .weight_en(weight_en));
SA22 U24_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_11_1), .partial_sum_in12(reg_psum23_11_2), .weight_in11(reg_weight23_11_1), .weight_in12(reg_weight23_11_2), .activation_in11(reg_activation24_10_1), .activation_in21(reg_activation24_10_2), .reg_partial_sum21(reg_psum24_11_1), .reg_partial_sum22(reg_psum24_11_2), .reg_weight21(reg_weight24_11_1), .reg_weight22(reg_weight24_11_2), .reg_activation12(reg_activation24_11_1), .reg_activation22(reg_activation24_11_2), .weight_en(weight_en));
SA22 U24_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_12_1), .partial_sum_in12(reg_psum23_12_2), .weight_in11(reg_weight23_12_1), .weight_in12(reg_weight23_12_2), .activation_in11(reg_activation24_11_1), .activation_in21(reg_activation24_11_2), .reg_partial_sum21(reg_psum24_12_1), .reg_partial_sum22(reg_psum24_12_2), .reg_weight21(reg_weight24_12_1), .reg_weight22(reg_weight24_12_2), .reg_activation12(reg_activation24_12_1), .reg_activation22(reg_activation24_12_2), .weight_en(weight_en));
SA22 U24_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_13_1), .partial_sum_in12(reg_psum23_13_2), .weight_in11(reg_weight23_13_1), .weight_in12(reg_weight23_13_2), .activation_in11(reg_activation24_12_1), .activation_in21(reg_activation24_12_2), .reg_partial_sum21(reg_psum24_13_1), .reg_partial_sum22(reg_psum24_13_2), .reg_weight21(reg_weight24_13_1), .reg_weight22(reg_weight24_13_2), .reg_activation12(reg_activation24_13_1), .reg_activation22(reg_activation24_13_2), .weight_en(weight_en));
SA22 U24_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_14_1), .partial_sum_in12(reg_psum23_14_2), .weight_in11(reg_weight23_14_1), .weight_in12(reg_weight23_14_2), .activation_in11(reg_activation24_13_1), .activation_in21(reg_activation24_13_2), .reg_partial_sum21(reg_psum24_14_1), .reg_partial_sum22(reg_psum24_14_2), .reg_weight21(reg_weight24_14_1), .reg_weight22(reg_weight24_14_2), .reg_activation12(reg_activation24_14_1), .reg_activation22(reg_activation24_14_2), .weight_en(weight_en));
SA22 U24_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_15_1), .partial_sum_in12(reg_psum23_15_2), .weight_in11(reg_weight23_15_1), .weight_in12(reg_weight23_15_2), .activation_in11(reg_activation24_14_1), .activation_in21(reg_activation24_14_2), .reg_partial_sum21(reg_psum24_15_1), .reg_partial_sum22(reg_psum24_15_2), .reg_weight21(reg_weight24_15_1), .reg_weight22(reg_weight24_15_2), .reg_activation12(reg_activation24_15_1), .reg_activation22(reg_activation24_15_2), .weight_en(weight_en));
SA22 U24_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_16_1), .partial_sum_in12(reg_psum23_16_2), .weight_in11(reg_weight23_16_1), .weight_in12(reg_weight23_16_2), .activation_in11(reg_activation24_15_1), .activation_in21(reg_activation24_15_2), .reg_partial_sum21(reg_psum24_16_1), .reg_partial_sum22(reg_psum24_16_2), .reg_weight21(reg_weight24_16_1), .reg_weight22(reg_weight24_16_2), .reg_activation12(reg_activation24_16_1), .reg_activation22(reg_activation24_16_2), .weight_en(weight_en));
SA22 U24_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_17_1), .partial_sum_in12(reg_psum23_17_2), .weight_in11(reg_weight23_17_1), .weight_in12(reg_weight23_17_2), .activation_in11(reg_activation24_16_1), .activation_in21(reg_activation24_16_2), .reg_partial_sum21(reg_psum24_17_1), .reg_partial_sum22(reg_psum24_17_2), .reg_weight21(reg_weight24_17_1), .reg_weight22(reg_weight24_17_2), .reg_activation12(reg_activation24_17_1), .reg_activation22(reg_activation24_17_2), .weight_en(weight_en));
SA22 U24_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_18_1), .partial_sum_in12(reg_psum23_18_2), .weight_in11(reg_weight23_18_1), .weight_in12(reg_weight23_18_2), .activation_in11(reg_activation24_17_1), .activation_in21(reg_activation24_17_2), .reg_partial_sum21(reg_psum24_18_1), .reg_partial_sum22(reg_psum24_18_2), .reg_weight21(reg_weight24_18_1), .reg_weight22(reg_weight24_18_2), .reg_activation12(reg_activation24_18_1), .reg_activation22(reg_activation24_18_2), .weight_en(weight_en));
SA22 U24_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_19_1), .partial_sum_in12(reg_psum23_19_2), .weight_in11(reg_weight23_19_1), .weight_in12(reg_weight23_19_2), .activation_in11(reg_activation24_18_1), .activation_in21(reg_activation24_18_2), .reg_partial_sum21(reg_psum24_19_1), .reg_partial_sum22(reg_psum24_19_2), .reg_weight21(reg_weight24_19_1), .reg_weight22(reg_weight24_19_2), .reg_activation12(reg_activation24_19_1), .reg_activation22(reg_activation24_19_2), .weight_en(weight_en));
SA22 U24_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_20_1), .partial_sum_in12(reg_psum23_20_2), .weight_in11(reg_weight23_20_1), .weight_in12(reg_weight23_20_2), .activation_in11(reg_activation24_19_1), .activation_in21(reg_activation24_19_2), .reg_partial_sum21(reg_psum24_20_1), .reg_partial_sum22(reg_psum24_20_2), .reg_weight21(reg_weight24_20_1), .reg_weight22(reg_weight24_20_2), .reg_activation12(reg_activation24_20_1), .reg_activation22(reg_activation24_20_2), .weight_en(weight_en));
SA22 U24_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_21_1), .partial_sum_in12(reg_psum23_21_2), .weight_in11(reg_weight23_21_1), .weight_in12(reg_weight23_21_2), .activation_in11(reg_activation24_20_1), .activation_in21(reg_activation24_20_2), .reg_partial_sum21(reg_psum24_21_1), .reg_partial_sum22(reg_psum24_21_2), .reg_weight21(reg_weight24_21_1), .reg_weight22(reg_weight24_21_2), .reg_activation12(reg_activation24_21_1), .reg_activation22(reg_activation24_21_2), .weight_en(weight_en));
SA22 U24_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_22_1), .partial_sum_in12(reg_psum23_22_2), .weight_in11(reg_weight23_22_1), .weight_in12(reg_weight23_22_2), .activation_in11(reg_activation24_21_1), .activation_in21(reg_activation24_21_2), .reg_partial_sum21(reg_psum24_22_1), .reg_partial_sum22(reg_psum24_22_2), .reg_weight21(reg_weight24_22_1), .reg_weight22(reg_weight24_22_2), .reg_activation12(reg_activation24_22_1), .reg_activation22(reg_activation24_22_2), .weight_en(weight_en));
SA22 U24_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_23_1), .partial_sum_in12(reg_psum23_23_2), .weight_in11(reg_weight23_23_1), .weight_in12(reg_weight23_23_2), .activation_in11(reg_activation24_22_1), .activation_in21(reg_activation24_22_2), .reg_partial_sum21(reg_psum24_23_1), .reg_partial_sum22(reg_psum24_23_2), .reg_weight21(reg_weight24_23_1), .reg_weight22(reg_weight24_23_2), .reg_activation12(reg_activation24_23_1), .reg_activation22(reg_activation24_23_2), .weight_en(weight_en));
SA22 U24_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_24_1), .partial_sum_in12(reg_psum23_24_2), .weight_in11(reg_weight23_24_1), .weight_in12(reg_weight23_24_2), .activation_in11(reg_activation24_23_1), .activation_in21(reg_activation24_23_2), .reg_partial_sum21(reg_psum24_24_1), .reg_partial_sum22(reg_psum24_24_2), .reg_weight21(reg_weight24_24_1), .reg_weight22(reg_weight24_24_2), .reg_activation12(reg_activation24_24_1), .reg_activation22(reg_activation24_24_2), .weight_en(weight_en));
SA22 U24_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_25_1), .partial_sum_in12(reg_psum23_25_2), .weight_in11(reg_weight23_25_1), .weight_in12(reg_weight23_25_2), .activation_in11(reg_activation24_24_1), .activation_in21(reg_activation24_24_2), .reg_partial_sum21(reg_psum24_25_1), .reg_partial_sum22(reg_psum24_25_2), .reg_weight21(reg_weight24_25_1), .reg_weight22(reg_weight24_25_2), .reg_activation12(reg_activation24_25_1), .reg_activation22(reg_activation24_25_2), .weight_en(weight_en));
SA22 U24_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_26_1), .partial_sum_in12(reg_psum23_26_2), .weight_in11(reg_weight23_26_1), .weight_in12(reg_weight23_26_2), .activation_in11(reg_activation24_25_1), .activation_in21(reg_activation24_25_2), .reg_partial_sum21(reg_psum24_26_1), .reg_partial_sum22(reg_psum24_26_2), .reg_weight21(reg_weight24_26_1), .reg_weight22(reg_weight24_26_2), .reg_activation12(reg_activation24_26_1), .reg_activation22(reg_activation24_26_2), .weight_en(weight_en));
SA22 U24_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_27_1), .partial_sum_in12(reg_psum23_27_2), .weight_in11(reg_weight23_27_1), .weight_in12(reg_weight23_27_2), .activation_in11(reg_activation24_26_1), .activation_in21(reg_activation24_26_2), .reg_partial_sum21(reg_psum24_27_1), .reg_partial_sum22(reg_psum24_27_2), .reg_weight21(reg_weight24_27_1), .reg_weight22(reg_weight24_27_2), .reg_activation12(reg_activation24_27_1), .reg_activation22(reg_activation24_27_2), .weight_en(weight_en));
SA22 U24_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_28_1), .partial_sum_in12(reg_psum23_28_2), .weight_in11(reg_weight23_28_1), .weight_in12(reg_weight23_28_2), .activation_in11(reg_activation24_27_1), .activation_in21(reg_activation24_27_2), .reg_partial_sum21(reg_psum24_28_1), .reg_partial_sum22(reg_psum24_28_2), .reg_weight21(reg_weight24_28_1), .reg_weight22(reg_weight24_28_2), .reg_activation12(reg_activation24_28_1), .reg_activation22(reg_activation24_28_2), .weight_en(weight_en));
SA22 U24_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_29_1), .partial_sum_in12(reg_psum23_29_2), .weight_in11(reg_weight23_29_1), .weight_in12(reg_weight23_29_2), .activation_in11(reg_activation24_28_1), .activation_in21(reg_activation24_28_2), .reg_partial_sum21(reg_psum24_29_1), .reg_partial_sum22(reg_psum24_29_2), .reg_weight21(reg_weight24_29_1), .reg_weight22(reg_weight24_29_2), .reg_activation12(reg_activation24_29_1), .reg_activation22(reg_activation24_29_2), .weight_en(weight_en));
SA22 U24_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_30_1), .partial_sum_in12(reg_psum23_30_2), .weight_in11(reg_weight23_30_1), .weight_in12(reg_weight23_30_2), .activation_in11(reg_activation24_29_1), .activation_in21(reg_activation24_29_2), .reg_partial_sum21(reg_psum24_30_1), .reg_partial_sum22(reg_psum24_30_2), .reg_weight21(reg_weight24_30_1), .reg_weight22(reg_weight24_30_2), .reg_activation12(reg_activation24_30_1), .reg_activation22(reg_activation24_30_2), .weight_en(weight_en));
SA22 U24_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_31_1), .partial_sum_in12(reg_psum23_31_2), .weight_in11(reg_weight23_31_1), .weight_in12(reg_weight23_31_2), .activation_in11(reg_activation24_30_1), .activation_in21(reg_activation24_30_2), .reg_partial_sum21(reg_psum24_31_1), .reg_partial_sum22(reg_psum24_31_2), .reg_weight21(reg_weight24_31_1), .reg_weight22(reg_weight24_31_2), .reg_activation12(reg_activation24_31_1), .reg_activation22(reg_activation24_31_2), .weight_en(weight_en));
SA22 U24_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum23_32_1), .partial_sum_in12(reg_psum23_32_2), .weight_in11(reg_weight23_32_1), .weight_in12(reg_weight23_32_2), .activation_in11(reg_activation24_31_1), .activation_in21(reg_activation24_31_2), .reg_partial_sum21(reg_psum24_32_1), .reg_partial_sum22(reg_psum24_32_2), .reg_weight21(reg_weight24_32_1), .reg_weight22(reg_weight24_32_2), .weight_en(weight_en));
SA22 U25_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_1_1), .partial_sum_in12(reg_psum24_1_2), .weight_in11(reg_weight24_1_1), .weight_in12(reg_weight24_1_2), .activation_in11(in_activation25_1_1), .activation_in21(in_activation25_1_2), .reg_partial_sum21(reg_psum25_1_1), .reg_partial_sum22(reg_psum25_1_2), .reg_weight21(reg_weight25_1_1), .reg_weight22(reg_weight25_1_2), .reg_activation12(reg_activation25_1_1), .reg_activation22(reg_activation25_1_2), .weight_en(weight_en));
SA22 U25_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_2_1), .partial_sum_in12(reg_psum24_2_2), .weight_in11(reg_weight24_2_1), .weight_in12(reg_weight24_2_2), .activation_in11(reg_activation25_1_1), .activation_in21(reg_activation25_1_2), .reg_partial_sum21(reg_psum25_2_1), .reg_partial_sum22(reg_psum25_2_2), .reg_weight21(reg_weight25_2_1), .reg_weight22(reg_weight25_2_2), .reg_activation12(reg_activation25_2_1), .reg_activation22(reg_activation25_2_2), .weight_en(weight_en));
SA22 U25_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_3_1), .partial_sum_in12(reg_psum24_3_2), .weight_in11(reg_weight24_3_1), .weight_in12(reg_weight24_3_2), .activation_in11(reg_activation25_2_1), .activation_in21(reg_activation25_2_2), .reg_partial_sum21(reg_psum25_3_1), .reg_partial_sum22(reg_psum25_3_2), .reg_weight21(reg_weight25_3_1), .reg_weight22(reg_weight25_3_2), .reg_activation12(reg_activation25_3_1), .reg_activation22(reg_activation25_3_2), .weight_en(weight_en));
SA22 U25_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_4_1), .partial_sum_in12(reg_psum24_4_2), .weight_in11(reg_weight24_4_1), .weight_in12(reg_weight24_4_2), .activation_in11(reg_activation25_3_1), .activation_in21(reg_activation25_3_2), .reg_partial_sum21(reg_psum25_4_1), .reg_partial_sum22(reg_psum25_4_2), .reg_weight21(reg_weight25_4_1), .reg_weight22(reg_weight25_4_2), .reg_activation12(reg_activation25_4_1), .reg_activation22(reg_activation25_4_2), .weight_en(weight_en));
SA22 U25_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_5_1), .partial_sum_in12(reg_psum24_5_2), .weight_in11(reg_weight24_5_1), .weight_in12(reg_weight24_5_2), .activation_in11(reg_activation25_4_1), .activation_in21(reg_activation25_4_2), .reg_partial_sum21(reg_psum25_5_1), .reg_partial_sum22(reg_psum25_5_2), .reg_weight21(reg_weight25_5_1), .reg_weight22(reg_weight25_5_2), .reg_activation12(reg_activation25_5_1), .reg_activation22(reg_activation25_5_2), .weight_en(weight_en));
SA22 U25_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_6_1), .partial_sum_in12(reg_psum24_6_2), .weight_in11(reg_weight24_6_1), .weight_in12(reg_weight24_6_2), .activation_in11(reg_activation25_5_1), .activation_in21(reg_activation25_5_2), .reg_partial_sum21(reg_psum25_6_1), .reg_partial_sum22(reg_psum25_6_2), .reg_weight21(reg_weight25_6_1), .reg_weight22(reg_weight25_6_2), .reg_activation12(reg_activation25_6_1), .reg_activation22(reg_activation25_6_2), .weight_en(weight_en));
SA22 U25_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_7_1), .partial_sum_in12(reg_psum24_7_2), .weight_in11(reg_weight24_7_1), .weight_in12(reg_weight24_7_2), .activation_in11(reg_activation25_6_1), .activation_in21(reg_activation25_6_2), .reg_partial_sum21(reg_psum25_7_1), .reg_partial_sum22(reg_psum25_7_2), .reg_weight21(reg_weight25_7_1), .reg_weight22(reg_weight25_7_2), .reg_activation12(reg_activation25_7_1), .reg_activation22(reg_activation25_7_2), .weight_en(weight_en));
SA22 U25_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_8_1), .partial_sum_in12(reg_psum24_8_2), .weight_in11(reg_weight24_8_1), .weight_in12(reg_weight24_8_2), .activation_in11(reg_activation25_7_1), .activation_in21(reg_activation25_7_2), .reg_partial_sum21(reg_psum25_8_1), .reg_partial_sum22(reg_psum25_8_2), .reg_weight21(reg_weight25_8_1), .reg_weight22(reg_weight25_8_2), .reg_activation12(reg_activation25_8_1), .reg_activation22(reg_activation25_8_2), .weight_en(weight_en));
SA22 U25_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_9_1), .partial_sum_in12(reg_psum24_9_2), .weight_in11(reg_weight24_9_1), .weight_in12(reg_weight24_9_2), .activation_in11(reg_activation25_8_1), .activation_in21(reg_activation25_8_2), .reg_partial_sum21(reg_psum25_9_1), .reg_partial_sum22(reg_psum25_9_2), .reg_weight21(reg_weight25_9_1), .reg_weight22(reg_weight25_9_2), .reg_activation12(reg_activation25_9_1), .reg_activation22(reg_activation25_9_2), .weight_en(weight_en));
SA22 U25_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_10_1), .partial_sum_in12(reg_psum24_10_2), .weight_in11(reg_weight24_10_1), .weight_in12(reg_weight24_10_2), .activation_in11(reg_activation25_9_1), .activation_in21(reg_activation25_9_2), .reg_partial_sum21(reg_psum25_10_1), .reg_partial_sum22(reg_psum25_10_2), .reg_weight21(reg_weight25_10_1), .reg_weight22(reg_weight25_10_2), .reg_activation12(reg_activation25_10_1), .reg_activation22(reg_activation25_10_2), .weight_en(weight_en));
SA22 U25_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_11_1), .partial_sum_in12(reg_psum24_11_2), .weight_in11(reg_weight24_11_1), .weight_in12(reg_weight24_11_2), .activation_in11(reg_activation25_10_1), .activation_in21(reg_activation25_10_2), .reg_partial_sum21(reg_psum25_11_1), .reg_partial_sum22(reg_psum25_11_2), .reg_weight21(reg_weight25_11_1), .reg_weight22(reg_weight25_11_2), .reg_activation12(reg_activation25_11_1), .reg_activation22(reg_activation25_11_2), .weight_en(weight_en));
SA22 U25_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_12_1), .partial_sum_in12(reg_psum24_12_2), .weight_in11(reg_weight24_12_1), .weight_in12(reg_weight24_12_2), .activation_in11(reg_activation25_11_1), .activation_in21(reg_activation25_11_2), .reg_partial_sum21(reg_psum25_12_1), .reg_partial_sum22(reg_psum25_12_2), .reg_weight21(reg_weight25_12_1), .reg_weight22(reg_weight25_12_2), .reg_activation12(reg_activation25_12_1), .reg_activation22(reg_activation25_12_2), .weight_en(weight_en));
SA22 U25_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_13_1), .partial_sum_in12(reg_psum24_13_2), .weight_in11(reg_weight24_13_1), .weight_in12(reg_weight24_13_2), .activation_in11(reg_activation25_12_1), .activation_in21(reg_activation25_12_2), .reg_partial_sum21(reg_psum25_13_1), .reg_partial_sum22(reg_psum25_13_2), .reg_weight21(reg_weight25_13_1), .reg_weight22(reg_weight25_13_2), .reg_activation12(reg_activation25_13_1), .reg_activation22(reg_activation25_13_2), .weight_en(weight_en));
SA22 U25_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_14_1), .partial_sum_in12(reg_psum24_14_2), .weight_in11(reg_weight24_14_1), .weight_in12(reg_weight24_14_2), .activation_in11(reg_activation25_13_1), .activation_in21(reg_activation25_13_2), .reg_partial_sum21(reg_psum25_14_1), .reg_partial_sum22(reg_psum25_14_2), .reg_weight21(reg_weight25_14_1), .reg_weight22(reg_weight25_14_2), .reg_activation12(reg_activation25_14_1), .reg_activation22(reg_activation25_14_2), .weight_en(weight_en));
SA22 U25_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_15_1), .partial_sum_in12(reg_psum24_15_2), .weight_in11(reg_weight24_15_1), .weight_in12(reg_weight24_15_2), .activation_in11(reg_activation25_14_1), .activation_in21(reg_activation25_14_2), .reg_partial_sum21(reg_psum25_15_1), .reg_partial_sum22(reg_psum25_15_2), .reg_weight21(reg_weight25_15_1), .reg_weight22(reg_weight25_15_2), .reg_activation12(reg_activation25_15_1), .reg_activation22(reg_activation25_15_2), .weight_en(weight_en));
SA22 U25_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_16_1), .partial_sum_in12(reg_psum24_16_2), .weight_in11(reg_weight24_16_1), .weight_in12(reg_weight24_16_2), .activation_in11(reg_activation25_15_1), .activation_in21(reg_activation25_15_2), .reg_partial_sum21(reg_psum25_16_1), .reg_partial_sum22(reg_psum25_16_2), .reg_weight21(reg_weight25_16_1), .reg_weight22(reg_weight25_16_2), .reg_activation12(reg_activation25_16_1), .reg_activation22(reg_activation25_16_2), .weight_en(weight_en));
SA22 U25_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_17_1), .partial_sum_in12(reg_psum24_17_2), .weight_in11(reg_weight24_17_1), .weight_in12(reg_weight24_17_2), .activation_in11(reg_activation25_16_1), .activation_in21(reg_activation25_16_2), .reg_partial_sum21(reg_psum25_17_1), .reg_partial_sum22(reg_psum25_17_2), .reg_weight21(reg_weight25_17_1), .reg_weight22(reg_weight25_17_2), .reg_activation12(reg_activation25_17_1), .reg_activation22(reg_activation25_17_2), .weight_en(weight_en));
SA22 U25_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_18_1), .partial_sum_in12(reg_psum24_18_2), .weight_in11(reg_weight24_18_1), .weight_in12(reg_weight24_18_2), .activation_in11(reg_activation25_17_1), .activation_in21(reg_activation25_17_2), .reg_partial_sum21(reg_psum25_18_1), .reg_partial_sum22(reg_psum25_18_2), .reg_weight21(reg_weight25_18_1), .reg_weight22(reg_weight25_18_2), .reg_activation12(reg_activation25_18_1), .reg_activation22(reg_activation25_18_2), .weight_en(weight_en));
SA22 U25_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_19_1), .partial_sum_in12(reg_psum24_19_2), .weight_in11(reg_weight24_19_1), .weight_in12(reg_weight24_19_2), .activation_in11(reg_activation25_18_1), .activation_in21(reg_activation25_18_2), .reg_partial_sum21(reg_psum25_19_1), .reg_partial_sum22(reg_psum25_19_2), .reg_weight21(reg_weight25_19_1), .reg_weight22(reg_weight25_19_2), .reg_activation12(reg_activation25_19_1), .reg_activation22(reg_activation25_19_2), .weight_en(weight_en));
SA22 U25_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_20_1), .partial_sum_in12(reg_psum24_20_2), .weight_in11(reg_weight24_20_1), .weight_in12(reg_weight24_20_2), .activation_in11(reg_activation25_19_1), .activation_in21(reg_activation25_19_2), .reg_partial_sum21(reg_psum25_20_1), .reg_partial_sum22(reg_psum25_20_2), .reg_weight21(reg_weight25_20_1), .reg_weight22(reg_weight25_20_2), .reg_activation12(reg_activation25_20_1), .reg_activation22(reg_activation25_20_2), .weight_en(weight_en));
SA22 U25_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_21_1), .partial_sum_in12(reg_psum24_21_2), .weight_in11(reg_weight24_21_1), .weight_in12(reg_weight24_21_2), .activation_in11(reg_activation25_20_1), .activation_in21(reg_activation25_20_2), .reg_partial_sum21(reg_psum25_21_1), .reg_partial_sum22(reg_psum25_21_2), .reg_weight21(reg_weight25_21_1), .reg_weight22(reg_weight25_21_2), .reg_activation12(reg_activation25_21_1), .reg_activation22(reg_activation25_21_2), .weight_en(weight_en));
SA22 U25_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_22_1), .partial_sum_in12(reg_psum24_22_2), .weight_in11(reg_weight24_22_1), .weight_in12(reg_weight24_22_2), .activation_in11(reg_activation25_21_1), .activation_in21(reg_activation25_21_2), .reg_partial_sum21(reg_psum25_22_1), .reg_partial_sum22(reg_psum25_22_2), .reg_weight21(reg_weight25_22_1), .reg_weight22(reg_weight25_22_2), .reg_activation12(reg_activation25_22_1), .reg_activation22(reg_activation25_22_2), .weight_en(weight_en));
SA22 U25_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_23_1), .partial_sum_in12(reg_psum24_23_2), .weight_in11(reg_weight24_23_1), .weight_in12(reg_weight24_23_2), .activation_in11(reg_activation25_22_1), .activation_in21(reg_activation25_22_2), .reg_partial_sum21(reg_psum25_23_1), .reg_partial_sum22(reg_psum25_23_2), .reg_weight21(reg_weight25_23_1), .reg_weight22(reg_weight25_23_2), .reg_activation12(reg_activation25_23_1), .reg_activation22(reg_activation25_23_2), .weight_en(weight_en));
SA22 U25_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_24_1), .partial_sum_in12(reg_psum24_24_2), .weight_in11(reg_weight24_24_1), .weight_in12(reg_weight24_24_2), .activation_in11(reg_activation25_23_1), .activation_in21(reg_activation25_23_2), .reg_partial_sum21(reg_psum25_24_1), .reg_partial_sum22(reg_psum25_24_2), .reg_weight21(reg_weight25_24_1), .reg_weight22(reg_weight25_24_2), .reg_activation12(reg_activation25_24_1), .reg_activation22(reg_activation25_24_2), .weight_en(weight_en));
SA22 U25_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_25_1), .partial_sum_in12(reg_psum24_25_2), .weight_in11(reg_weight24_25_1), .weight_in12(reg_weight24_25_2), .activation_in11(reg_activation25_24_1), .activation_in21(reg_activation25_24_2), .reg_partial_sum21(reg_psum25_25_1), .reg_partial_sum22(reg_psum25_25_2), .reg_weight21(reg_weight25_25_1), .reg_weight22(reg_weight25_25_2), .reg_activation12(reg_activation25_25_1), .reg_activation22(reg_activation25_25_2), .weight_en(weight_en));
SA22 U25_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_26_1), .partial_sum_in12(reg_psum24_26_2), .weight_in11(reg_weight24_26_1), .weight_in12(reg_weight24_26_2), .activation_in11(reg_activation25_25_1), .activation_in21(reg_activation25_25_2), .reg_partial_sum21(reg_psum25_26_1), .reg_partial_sum22(reg_psum25_26_2), .reg_weight21(reg_weight25_26_1), .reg_weight22(reg_weight25_26_2), .reg_activation12(reg_activation25_26_1), .reg_activation22(reg_activation25_26_2), .weight_en(weight_en));
SA22 U25_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_27_1), .partial_sum_in12(reg_psum24_27_2), .weight_in11(reg_weight24_27_1), .weight_in12(reg_weight24_27_2), .activation_in11(reg_activation25_26_1), .activation_in21(reg_activation25_26_2), .reg_partial_sum21(reg_psum25_27_1), .reg_partial_sum22(reg_psum25_27_2), .reg_weight21(reg_weight25_27_1), .reg_weight22(reg_weight25_27_2), .reg_activation12(reg_activation25_27_1), .reg_activation22(reg_activation25_27_2), .weight_en(weight_en));
SA22 U25_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_28_1), .partial_sum_in12(reg_psum24_28_2), .weight_in11(reg_weight24_28_1), .weight_in12(reg_weight24_28_2), .activation_in11(reg_activation25_27_1), .activation_in21(reg_activation25_27_2), .reg_partial_sum21(reg_psum25_28_1), .reg_partial_sum22(reg_psum25_28_2), .reg_weight21(reg_weight25_28_1), .reg_weight22(reg_weight25_28_2), .reg_activation12(reg_activation25_28_1), .reg_activation22(reg_activation25_28_2), .weight_en(weight_en));
SA22 U25_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_29_1), .partial_sum_in12(reg_psum24_29_2), .weight_in11(reg_weight24_29_1), .weight_in12(reg_weight24_29_2), .activation_in11(reg_activation25_28_1), .activation_in21(reg_activation25_28_2), .reg_partial_sum21(reg_psum25_29_1), .reg_partial_sum22(reg_psum25_29_2), .reg_weight21(reg_weight25_29_1), .reg_weight22(reg_weight25_29_2), .reg_activation12(reg_activation25_29_1), .reg_activation22(reg_activation25_29_2), .weight_en(weight_en));
SA22 U25_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_30_1), .partial_sum_in12(reg_psum24_30_2), .weight_in11(reg_weight24_30_1), .weight_in12(reg_weight24_30_2), .activation_in11(reg_activation25_29_1), .activation_in21(reg_activation25_29_2), .reg_partial_sum21(reg_psum25_30_1), .reg_partial_sum22(reg_psum25_30_2), .reg_weight21(reg_weight25_30_1), .reg_weight22(reg_weight25_30_2), .reg_activation12(reg_activation25_30_1), .reg_activation22(reg_activation25_30_2), .weight_en(weight_en));
SA22 U25_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_31_1), .partial_sum_in12(reg_psum24_31_2), .weight_in11(reg_weight24_31_1), .weight_in12(reg_weight24_31_2), .activation_in11(reg_activation25_30_1), .activation_in21(reg_activation25_30_2), .reg_partial_sum21(reg_psum25_31_1), .reg_partial_sum22(reg_psum25_31_2), .reg_weight21(reg_weight25_31_1), .reg_weight22(reg_weight25_31_2), .reg_activation12(reg_activation25_31_1), .reg_activation22(reg_activation25_31_2), .weight_en(weight_en));
SA22 U25_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum24_32_1), .partial_sum_in12(reg_psum24_32_2), .weight_in11(reg_weight24_32_1), .weight_in12(reg_weight24_32_2), .activation_in11(reg_activation25_31_1), .activation_in21(reg_activation25_31_2), .reg_partial_sum21(reg_psum25_32_1), .reg_partial_sum22(reg_psum25_32_2), .reg_weight21(reg_weight25_32_1), .reg_weight22(reg_weight25_32_2), .weight_en(weight_en));
SA22 U26_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_1_1), .partial_sum_in12(reg_psum25_1_2), .weight_in11(reg_weight25_1_1), .weight_in12(reg_weight25_1_2), .activation_in11(in_activation26_1_1), .activation_in21(in_activation26_1_2), .reg_partial_sum21(reg_psum26_1_1), .reg_partial_sum22(reg_psum26_1_2), .reg_weight21(reg_weight26_1_1), .reg_weight22(reg_weight26_1_2), .reg_activation12(reg_activation26_1_1), .reg_activation22(reg_activation26_1_2), .weight_en(weight_en));
SA22 U26_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_2_1), .partial_sum_in12(reg_psum25_2_2), .weight_in11(reg_weight25_2_1), .weight_in12(reg_weight25_2_2), .activation_in11(reg_activation26_1_1), .activation_in21(reg_activation26_1_2), .reg_partial_sum21(reg_psum26_2_1), .reg_partial_sum22(reg_psum26_2_2), .reg_weight21(reg_weight26_2_1), .reg_weight22(reg_weight26_2_2), .reg_activation12(reg_activation26_2_1), .reg_activation22(reg_activation26_2_2), .weight_en(weight_en));
SA22 U26_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_3_1), .partial_sum_in12(reg_psum25_3_2), .weight_in11(reg_weight25_3_1), .weight_in12(reg_weight25_3_2), .activation_in11(reg_activation26_2_1), .activation_in21(reg_activation26_2_2), .reg_partial_sum21(reg_psum26_3_1), .reg_partial_sum22(reg_psum26_3_2), .reg_weight21(reg_weight26_3_1), .reg_weight22(reg_weight26_3_2), .reg_activation12(reg_activation26_3_1), .reg_activation22(reg_activation26_3_2), .weight_en(weight_en));
SA22 U26_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_4_1), .partial_sum_in12(reg_psum25_4_2), .weight_in11(reg_weight25_4_1), .weight_in12(reg_weight25_4_2), .activation_in11(reg_activation26_3_1), .activation_in21(reg_activation26_3_2), .reg_partial_sum21(reg_psum26_4_1), .reg_partial_sum22(reg_psum26_4_2), .reg_weight21(reg_weight26_4_1), .reg_weight22(reg_weight26_4_2), .reg_activation12(reg_activation26_4_1), .reg_activation22(reg_activation26_4_2), .weight_en(weight_en));
SA22 U26_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_5_1), .partial_sum_in12(reg_psum25_5_2), .weight_in11(reg_weight25_5_1), .weight_in12(reg_weight25_5_2), .activation_in11(reg_activation26_4_1), .activation_in21(reg_activation26_4_2), .reg_partial_sum21(reg_psum26_5_1), .reg_partial_sum22(reg_psum26_5_2), .reg_weight21(reg_weight26_5_1), .reg_weight22(reg_weight26_5_2), .reg_activation12(reg_activation26_5_1), .reg_activation22(reg_activation26_5_2), .weight_en(weight_en));
SA22 U26_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_6_1), .partial_sum_in12(reg_psum25_6_2), .weight_in11(reg_weight25_6_1), .weight_in12(reg_weight25_6_2), .activation_in11(reg_activation26_5_1), .activation_in21(reg_activation26_5_2), .reg_partial_sum21(reg_psum26_6_1), .reg_partial_sum22(reg_psum26_6_2), .reg_weight21(reg_weight26_6_1), .reg_weight22(reg_weight26_6_2), .reg_activation12(reg_activation26_6_1), .reg_activation22(reg_activation26_6_2), .weight_en(weight_en));
SA22 U26_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_7_1), .partial_sum_in12(reg_psum25_7_2), .weight_in11(reg_weight25_7_1), .weight_in12(reg_weight25_7_2), .activation_in11(reg_activation26_6_1), .activation_in21(reg_activation26_6_2), .reg_partial_sum21(reg_psum26_7_1), .reg_partial_sum22(reg_psum26_7_2), .reg_weight21(reg_weight26_7_1), .reg_weight22(reg_weight26_7_2), .reg_activation12(reg_activation26_7_1), .reg_activation22(reg_activation26_7_2), .weight_en(weight_en));
SA22 U26_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_8_1), .partial_sum_in12(reg_psum25_8_2), .weight_in11(reg_weight25_8_1), .weight_in12(reg_weight25_8_2), .activation_in11(reg_activation26_7_1), .activation_in21(reg_activation26_7_2), .reg_partial_sum21(reg_psum26_8_1), .reg_partial_sum22(reg_psum26_8_2), .reg_weight21(reg_weight26_8_1), .reg_weight22(reg_weight26_8_2), .reg_activation12(reg_activation26_8_1), .reg_activation22(reg_activation26_8_2), .weight_en(weight_en));
SA22 U26_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_9_1), .partial_sum_in12(reg_psum25_9_2), .weight_in11(reg_weight25_9_1), .weight_in12(reg_weight25_9_2), .activation_in11(reg_activation26_8_1), .activation_in21(reg_activation26_8_2), .reg_partial_sum21(reg_psum26_9_1), .reg_partial_sum22(reg_psum26_9_2), .reg_weight21(reg_weight26_9_1), .reg_weight22(reg_weight26_9_2), .reg_activation12(reg_activation26_9_1), .reg_activation22(reg_activation26_9_2), .weight_en(weight_en));
SA22 U26_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_10_1), .partial_sum_in12(reg_psum25_10_2), .weight_in11(reg_weight25_10_1), .weight_in12(reg_weight25_10_2), .activation_in11(reg_activation26_9_1), .activation_in21(reg_activation26_9_2), .reg_partial_sum21(reg_psum26_10_1), .reg_partial_sum22(reg_psum26_10_2), .reg_weight21(reg_weight26_10_1), .reg_weight22(reg_weight26_10_2), .reg_activation12(reg_activation26_10_1), .reg_activation22(reg_activation26_10_2), .weight_en(weight_en));
SA22 U26_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_11_1), .partial_sum_in12(reg_psum25_11_2), .weight_in11(reg_weight25_11_1), .weight_in12(reg_weight25_11_2), .activation_in11(reg_activation26_10_1), .activation_in21(reg_activation26_10_2), .reg_partial_sum21(reg_psum26_11_1), .reg_partial_sum22(reg_psum26_11_2), .reg_weight21(reg_weight26_11_1), .reg_weight22(reg_weight26_11_2), .reg_activation12(reg_activation26_11_1), .reg_activation22(reg_activation26_11_2), .weight_en(weight_en));
SA22 U26_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_12_1), .partial_sum_in12(reg_psum25_12_2), .weight_in11(reg_weight25_12_1), .weight_in12(reg_weight25_12_2), .activation_in11(reg_activation26_11_1), .activation_in21(reg_activation26_11_2), .reg_partial_sum21(reg_psum26_12_1), .reg_partial_sum22(reg_psum26_12_2), .reg_weight21(reg_weight26_12_1), .reg_weight22(reg_weight26_12_2), .reg_activation12(reg_activation26_12_1), .reg_activation22(reg_activation26_12_2), .weight_en(weight_en));
SA22 U26_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_13_1), .partial_sum_in12(reg_psum25_13_2), .weight_in11(reg_weight25_13_1), .weight_in12(reg_weight25_13_2), .activation_in11(reg_activation26_12_1), .activation_in21(reg_activation26_12_2), .reg_partial_sum21(reg_psum26_13_1), .reg_partial_sum22(reg_psum26_13_2), .reg_weight21(reg_weight26_13_1), .reg_weight22(reg_weight26_13_2), .reg_activation12(reg_activation26_13_1), .reg_activation22(reg_activation26_13_2), .weight_en(weight_en));
SA22 U26_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_14_1), .partial_sum_in12(reg_psum25_14_2), .weight_in11(reg_weight25_14_1), .weight_in12(reg_weight25_14_2), .activation_in11(reg_activation26_13_1), .activation_in21(reg_activation26_13_2), .reg_partial_sum21(reg_psum26_14_1), .reg_partial_sum22(reg_psum26_14_2), .reg_weight21(reg_weight26_14_1), .reg_weight22(reg_weight26_14_2), .reg_activation12(reg_activation26_14_1), .reg_activation22(reg_activation26_14_2), .weight_en(weight_en));
SA22 U26_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_15_1), .partial_sum_in12(reg_psum25_15_2), .weight_in11(reg_weight25_15_1), .weight_in12(reg_weight25_15_2), .activation_in11(reg_activation26_14_1), .activation_in21(reg_activation26_14_2), .reg_partial_sum21(reg_psum26_15_1), .reg_partial_sum22(reg_psum26_15_2), .reg_weight21(reg_weight26_15_1), .reg_weight22(reg_weight26_15_2), .reg_activation12(reg_activation26_15_1), .reg_activation22(reg_activation26_15_2), .weight_en(weight_en));
SA22 U26_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_16_1), .partial_sum_in12(reg_psum25_16_2), .weight_in11(reg_weight25_16_1), .weight_in12(reg_weight25_16_2), .activation_in11(reg_activation26_15_1), .activation_in21(reg_activation26_15_2), .reg_partial_sum21(reg_psum26_16_1), .reg_partial_sum22(reg_psum26_16_2), .reg_weight21(reg_weight26_16_1), .reg_weight22(reg_weight26_16_2), .reg_activation12(reg_activation26_16_1), .reg_activation22(reg_activation26_16_2), .weight_en(weight_en));
SA22 U26_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_17_1), .partial_sum_in12(reg_psum25_17_2), .weight_in11(reg_weight25_17_1), .weight_in12(reg_weight25_17_2), .activation_in11(reg_activation26_16_1), .activation_in21(reg_activation26_16_2), .reg_partial_sum21(reg_psum26_17_1), .reg_partial_sum22(reg_psum26_17_2), .reg_weight21(reg_weight26_17_1), .reg_weight22(reg_weight26_17_2), .reg_activation12(reg_activation26_17_1), .reg_activation22(reg_activation26_17_2), .weight_en(weight_en));
SA22 U26_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_18_1), .partial_sum_in12(reg_psum25_18_2), .weight_in11(reg_weight25_18_1), .weight_in12(reg_weight25_18_2), .activation_in11(reg_activation26_17_1), .activation_in21(reg_activation26_17_2), .reg_partial_sum21(reg_psum26_18_1), .reg_partial_sum22(reg_psum26_18_2), .reg_weight21(reg_weight26_18_1), .reg_weight22(reg_weight26_18_2), .reg_activation12(reg_activation26_18_1), .reg_activation22(reg_activation26_18_2), .weight_en(weight_en));
SA22 U26_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_19_1), .partial_sum_in12(reg_psum25_19_2), .weight_in11(reg_weight25_19_1), .weight_in12(reg_weight25_19_2), .activation_in11(reg_activation26_18_1), .activation_in21(reg_activation26_18_2), .reg_partial_sum21(reg_psum26_19_1), .reg_partial_sum22(reg_psum26_19_2), .reg_weight21(reg_weight26_19_1), .reg_weight22(reg_weight26_19_2), .reg_activation12(reg_activation26_19_1), .reg_activation22(reg_activation26_19_2), .weight_en(weight_en));
SA22 U26_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_20_1), .partial_sum_in12(reg_psum25_20_2), .weight_in11(reg_weight25_20_1), .weight_in12(reg_weight25_20_2), .activation_in11(reg_activation26_19_1), .activation_in21(reg_activation26_19_2), .reg_partial_sum21(reg_psum26_20_1), .reg_partial_sum22(reg_psum26_20_2), .reg_weight21(reg_weight26_20_1), .reg_weight22(reg_weight26_20_2), .reg_activation12(reg_activation26_20_1), .reg_activation22(reg_activation26_20_2), .weight_en(weight_en));
SA22 U26_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_21_1), .partial_sum_in12(reg_psum25_21_2), .weight_in11(reg_weight25_21_1), .weight_in12(reg_weight25_21_2), .activation_in11(reg_activation26_20_1), .activation_in21(reg_activation26_20_2), .reg_partial_sum21(reg_psum26_21_1), .reg_partial_sum22(reg_psum26_21_2), .reg_weight21(reg_weight26_21_1), .reg_weight22(reg_weight26_21_2), .reg_activation12(reg_activation26_21_1), .reg_activation22(reg_activation26_21_2), .weight_en(weight_en));
SA22 U26_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_22_1), .partial_sum_in12(reg_psum25_22_2), .weight_in11(reg_weight25_22_1), .weight_in12(reg_weight25_22_2), .activation_in11(reg_activation26_21_1), .activation_in21(reg_activation26_21_2), .reg_partial_sum21(reg_psum26_22_1), .reg_partial_sum22(reg_psum26_22_2), .reg_weight21(reg_weight26_22_1), .reg_weight22(reg_weight26_22_2), .reg_activation12(reg_activation26_22_1), .reg_activation22(reg_activation26_22_2), .weight_en(weight_en));
SA22 U26_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_23_1), .partial_sum_in12(reg_psum25_23_2), .weight_in11(reg_weight25_23_1), .weight_in12(reg_weight25_23_2), .activation_in11(reg_activation26_22_1), .activation_in21(reg_activation26_22_2), .reg_partial_sum21(reg_psum26_23_1), .reg_partial_sum22(reg_psum26_23_2), .reg_weight21(reg_weight26_23_1), .reg_weight22(reg_weight26_23_2), .reg_activation12(reg_activation26_23_1), .reg_activation22(reg_activation26_23_2), .weight_en(weight_en));
SA22 U26_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_24_1), .partial_sum_in12(reg_psum25_24_2), .weight_in11(reg_weight25_24_1), .weight_in12(reg_weight25_24_2), .activation_in11(reg_activation26_23_1), .activation_in21(reg_activation26_23_2), .reg_partial_sum21(reg_psum26_24_1), .reg_partial_sum22(reg_psum26_24_2), .reg_weight21(reg_weight26_24_1), .reg_weight22(reg_weight26_24_2), .reg_activation12(reg_activation26_24_1), .reg_activation22(reg_activation26_24_2), .weight_en(weight_en));
SA22 U26_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_25_1), .partial_sum_in12(reg_psum25_25_2), .weight_in11(reg_weight25_25_1), .weight_in12(reg_weight25_25_2), .activation_in11(reg_activation26_24_1), .activation_in21(reg_activation26_24_2), .reg_partial_sum21(reg_psum26_25_1), .reg_partial_sum22(reg_psum26_25_2), .reg_weight21(reg_weight26_25_1), .reg_weight22(reg_weight26_25_2), .reg_activation12(reg_activation26_25_1), .reg_activation22(reg_activation26_25_2), .weight_en(weight_en));
SA22 U26_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_26_1), .partial_sum_in12(reg_psum25_26_2), .weight_in11(reg_weight25_26_1), .weight_in12(reg_weight25_26_2), .activation_in11(reg_activation26_25_1), .activation_in21(reg_activation26_25_2), .reg_partial_sum21(reg_psum26_26_1), .reg_partial_sum22(reg_psum26_26_2), .reg_weight21(reg_weight26_26_1), .reg_weight22(reg_weight26_26_2), .reg_activation12(reg_activation26_26_1), .reg_activation22(reg_activation26_26_2), .weight_en(weight_en));
SA22 U26_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_27_1), .partial_sum_in12(reg_psum25_27_2), .weight_in11(reg_weight25_27_1), .weight_in12(reg_weight25_27_2), .activation_in11(reg_activation26_26_1), .activation_in21(reg_activation26_26_2), .reg_partial_sum21(reg_psum26_27_1), .reg_partial_sum22(reg_psum26_27_2), .reg_weight21(reg_weight26_27_1), .reg_weight22(reg_weight26_27_2), .reg_activation12(reg_activation26_27_1), .reg_activation22(reg_activation26_27_2), .weight_en(weight_en));
SA22 U26_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_28_1), .partial_sum_in12(reg_psum25_28_2), .weight_in11(reg_weight25_28_1), .weight_in12(reg_weight25_28_2), .activation_in11(reg_activation26_27_1), .activation_in21(reg_activation26_27_2), .reg_partial_sum21(reg_psum26_28_1), .reg_partial_sum22(reg_psum26_28_2), .reg_weight21(reg_weight26_28_1), .reg_weight22(reg_weight26_28_2), .reg_activation12(reg_activation26_28_1), .reg_activation22(reg_activation26_28_2), .weight_en(weight_en));
SA22 U26_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_29_1), .partial_sum_in12(reg_psum25_29_2), .weight_in11(reg_weight25_29_1), .weight_in12(reg_weight25_29_2), .activation_in11(reg_activation26_28_1), .activation_in21(reg_activation26_28_2), .reg_partial_sum21(reg_psum26_29_1), .reg_partial_sum22(reg_psum26_29_2), .reg_weight21(reg_weight26_29_1), .reg_weight22(reg_weight26_29_2), .reg_activation12(reg_activation26_29_1), .reg_activation22(reg_activation26_29_2), .weight_en(weight_en));
SA22 U26_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_30_1), .partial_sum_in12(reg_psum25_30_2), .weight_in11(reg_weight25_30_1), .weight_in12(reg_weight25_30_2), .activation_in11(reg_activation26_29_1), .activation_in21(reg_activation26_29_2), .reg_partial_sum21(reg_psum26_30_1), .reg_partial_sum22(reg_psum26_30_2), .reg_weight21(reg_weight26_30_1), .reg_weight22(reg_weight26_30_2), .reg_activation12(reg_activation26_30_1), .reg_activation22(reg_activation26_30_2), .weight_en(weight_en));
SA22 U26_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_31_1), .partial_sum_in12(reg_psum25_31_2), .weight_in11(reg_weight25_31_1), .weight_in12(reg_weight25_31_2), .activation_in11(reg_activation26_30_1), .activation_in21(reg_activation26_30_2), .reg_partial_sum21(reg_psum26_31_1), .reg_partial_sum22(reg_psum26_31_2), .reg_weight21(reg_weight26_31_1), .reg_weight22(reg_weight26_31_2), .reg_activation12(reg_activation26_31_1), .reg_activation22(reg_activation26_31_2), .weight_en(weight_en));
SA22 U26_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum25_32_1), .partial_sum_in12(reg_psum25_32_2), .weight_in11(reg_weight25_32_1), .weight_in12(reg_weight25_32_2), .activation_in11(reg_activation26_31_1), .activation_in21(reg_activation26_31_2), .reg_partial_sum21(reg_psum26_32_1), .reg_partial_sum22(reg_psum26_32_2), .reg_weight21(reg_weight26_32_1), .reg_weight22(reg_weight26_32_2), .weight_en(weight_en));
SA22 U27_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_1_1), .partial_sum_in12(reg_psum26_1_2), .weight_in11(reg_weight26_1_1), .weight_in12(reg_weight26_1_2), .activation_in11(in_activation27_1_1), .activation_in21(in_activation27_1_2), .reg_partial_sum21(reg_psum27_1_1), .reg_partial_sum22(reg_psum27_1_2), .reg_weight21(reg_weight27_1_1), .reg_weight22(reg_weight27_1_2), .reg_activation12(reg_activation27_1_1), .reg_activation22(reg_activation27_1_2), .weight_en(weight_en));
SA22 U27_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_2_1), .partial_sum_in12(reg_psum26_2_2), .weight_in11(reg_weight26_2_1), .weight_in12(reg_weight26_2_2), .activation_in11(reg_activation27_1_1), .activation_in21(reg_activation27_1_2), .reg_partial_sum21(reg_psum27_2_1), .reg_partial_sum22(reg_psum27_2_2), .reg_weight21(reg_weight27_2_1), .reg_weight22(reg_weight27_2_2), .reg_activation12(reg_activation27_2_1), .reg_activation22(reg_activation27_2_2), .weight_en(weight_en));
SA22 U27_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_3_1), .partial_sum_in12(reg_psum26_3_2), .weight_in11(reg_weight26_3_1), .weight_in12(reg_weight26_3_2), .activation_in11(reg_activation27_2_1), .activation_in21(reg_activation27_2_2), .reg_partial_sum21(reg_psum27_3_1), .reg_partial_sum22(reg_psum27_3_2), .reg_weight21(reg_weight27_3_1), .reg_weight22(reg_weight27_3_2), .reg_activation12(reg_activation27_3_1), .reg_activation22(reg_activation27_3_2), .weight_en(weight_en));
SA22 U27_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_4_1), .partial_sum_in12(reg_psum26_4_2), .weight_in11(reg_weight26_4_1), .weight_in12(reg_weight26_4_2), .activation_in11(reg_activation27_3_1), .activation_in21(reg_activation27_3_2), .reg_partial_sum21(reg_psum27_4_1), .reg_partial_sum22(reg_psum27_4_2), .reg_weight21(reg_weight27_4_1), .reg_weight22(reg_weight27_4_2), .reg_activation12(reg_activation27_4_1), .reg_activation22(reg_activation27_4_2), .weight_en(weight_en));
SA22 U27_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_5_1), .partial_sum_in12(reg_psum26_5_2), .weight_in11(reg_weight26_5_1), .weight_in12(reg_weight26_5_2), .activation_in11(reg_activation27_4_1), .activation_in21(reg_activation27_4_2), .reg_partial_sum21(reg_psum27_5_1), .reg_partial_sum22(reg_psum27_5_2), .reg_weight21(reg_weight27_5_1), .reg_weight22(reg_weight27_5_2), .reg_activation12(reg_activation27_5_1), .reg_activation22(reg_activation27_5_2), .weight_en(weight_en));
SA22 U27_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_6_1), .partial_sum_in12(reg_psum26_6_2), .weight_in11(reg_weight26_6_1), .weight_in12(reg_weight26_6_2), .activation_in11(reg_activation27_5_1), .activation_in21(reg_activation27_5_2), .reg_partial_sum21(reg_psum27_6_1), .reg_partial_sum22(reg_psum27_6_2), .reg_weight21(reg_weight27_6_1), .reg_weight22(reg_weight27_6_2), .reg_activation12(reg_activation27_6_1), .reg_activation22(reg_activation27_6_2), .weight_en(weight_en));
SA22 U27_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_7_1), .partial_sum_in12(reg_psum26_7_2), .weight_in11(reg_weight26_7_1), .weight_in12(reg_weight26_7_2), .activation_in11(reg_activation27_6_1), .activation_in21(reg_activation27_6_2), .reg_partial_sum21(reg_psum27_7_1), .reg_partial_sum22(reg_psum27_7_2), .reg_weight21(reg_weight27_7_1), .reg_weight22(reg_weight27_7_2), .reg_activation12(reg_activation27_7_1), .reg_activation22(reg_activation27_7_2), .weight_en(weight_en));
SA22 U27_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_8_1), .partial_sum_in12(reg_psum26_8_2), .weight_in11(reg_weight26_8_1), .weight_in12(reg_weight26_8_2), .activation_in11(reg_activation27_7_1), .activation_in21(reg_activation27_7_2), .reg_partial_sum21(reg_psum27_8_1), .reg_partial_sum22(reg_psum27_8_2), .reg_weight21(reg_weight27_8_1), .reg_weight22(reg_weight27_8_2), .reg_activation12(reg_activation27_8_1), .reg_activation22(reg_activation27_8_2), .weight_en(weight_en));
SA22 U27_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_9_1), .partial_sum_in12(reg_psum26_9_2), .weight_in11(reg_weight26_9_1), .weight_in12(reg_weight26_9_2), .activation_in11(reg_activation27_8_1), .activation_in21(reg_activation27_8_2), .reg_partial_sum21(reg_psum27_9_1), .reg_partial_sum22(reg_psum27_9_2), .reg_weight21(reg_weight27_9_1), .reg_weight22(reg_weight27_9_2), .reg_activation12(reg_activation27_9_1), .reg_activation22(reg_activation27_9_2), .weight_en(weight_en));
SA22 U27_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_10_1), .partial_sum_in12(reg_psum26_10_2), .weight_in11(reg_weight26_10_1), .weight_in12(reg_weight26_10_2), .activation_in11(reg_activation27_9_1), .activation_in21(reg_activation27_9_2), .reg_partial_sum21(reg_psum27_10_1), .reg_partial_sum22(reg_psum27_10_2), .reg_weight21(reg_weight27_10_1), .reg_weight22(reg_weight27_10_2), .reg_activation12(reg_activation27_10_1), .reg_activation22(reg_activation27_10_2), .weight_en(weight_en));
SA22 U27_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_11_1), .partial_sum_in12(reg_psum26_11_2), .weight_in11(reg_weight26_11_1), .weight_in12(reg_weight26_11_2), .activation_in11(reg_activation27_10_1), .activation_in21(reg_activation27_10_2), .reg_partial_sum21(reg_psum27_11_1), .reg_partial_sum22(reg_psum27_11_2), .reg_weight21(reg_weight27_11_1), .reg_weight22(reg_weight27_11_2), .reg_activation12(reg_activation27_11_1), .reg_activation22(reg_activation27_11_2), .weight_en(weight_en));
SA22 U27_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_12_1), .partial_sum_in12(reg_psum26_12_2), .weight_in11(reg_weight26_12_1), .weight_in12(reg_weight26_12_2), .activation_in11(reg_activation27_11_1), .activation_in21(reg_activation27_11_2), .reg_partial_sum21(reg_psum27_12_1), .reg_partial_sum22(reg_psum27_12_2), .reg_weight21(reg_weight27_12_1), .reg_weight22(reg_weight27_12_2), .reg_activation12(reg_activation27_12_1), .reg_activation22(reg_activation27_12_2), .weight_en(weight_en));
SA22 U27_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_13_1), .partial_sum_in12(reg_psum26_13_2), .weight_in11(reg_weight26_13_1), .weight_in12(reg_weight26_13_2), .activation_in11(reg_activation27_12_1), .activation_in21(reg_activation27_12_2), .reg_partial_sum21(reg_psum27_13_1), .reg_partial_sum22(reg_psum27_13_2), .reg_weight21(reg_weight27_13_1), .reg_weight22(reg_weight27_13_2), .reg_activation12(reg_activation27_13_1), .reg_activation22(reg_activation27_13_2), .weight_en(weight_en));
SA22 U27_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_14_1), .partial_sum_in12(reg_psum26_14_2), .weight_in11(reg_weight26_14_1), .weight_in12(reg_weight26_14_2), .activation_in11(reg_activation27_13_1), .activation_in21(reg_activation27_13_2), .reg_partial_sum21(reg_psum27_14_1), .reg_partial_sum22(reg_psum27_14_2), .reg_weight21(reg_weight27_14_1), .reg_weight22(reg_weight27_14_2), .reg_activation12(reg_activation27_14_1), .reg_activation22(reg_activation27_14_2), .weight_en(weight_en));
SA22 U27_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_15_1), .partial_sum_in12(reg_psum26_15_2), .weight_in11(reg_weight26_15_1), .weight_in12(reg_weight26_15_2), .activation_in11(reg_activation27_14_1), .activation_in21(reg_activation27_14_2), .reg_partial_sum21(reg_psum27_15_1), .reg_partial_sum22(reg_psum27_15_2), .reg_weight21(reg_weight27_15_1), .reg_weight22(reg_weight27_15_2), .reg_activation12(reg_activation27_15_1), .reg_activation22(reg_activation27_15_2), .weight_en(weight_en));
SA22 U27_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_16_1), .partial_sum_in12(reg_psum26_16_2), .weight_in11(reg_weight26_16_1), .weight_in12(reg_weight26_16_2), .activation_in11(reg_activation27_15_1), .activation_in21(reg_activation27_15_2), .reg_partial_sum21(reg_psum27_16_1), .reg_partial_sum22(reg_psum27_16_2), .reg_weight21(reg_weight27_16_1), .reg_weight22(reg_weight27_16_2), .reg_activation12(reg_activation27_16_1), .reg_activation22(reg_activation27_16_2), .weight_en(weight_en));
SA22 U27_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_17_1), .partial_sum_in12(reg_psum26_17_2), .weight_in11(reg_weight26_17_1), .weight_in12(reg_weight26_17_2), .activation_in11(reg_activation27_16_1), .activation_in21(reg_activation27_16_2), .reg_partial_sum21(reg_psum27_17_1), .reg_partial_sum22(reg_psum27_17_2), .reg_weight21(reg_weight27_17_1), .reg_weight22(reg_weight27_17_2), .reg_activation12(reg_activation27_17_1), .reg_activation22(reg_activation27_17_2), .weight_en(weight_en));
SA22 U27_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_18_1), .partial_sum_in12(reg_psum26_18_2), .weight_in11(reg_weight26_18_1), .weight_in12(reg_weight26_18_2), .activation_in11(reg_activation27_17_1), .activation_in21(reg_activation27_17_2), .reg_partial_sum21(reg_psum27_18_1), .reg_partial_sum22(reg_psum27_18_2), .reg_weight21(reg_weight27_18_1), .reg_weight22(reg_weight27_18_2), .reg_activation12(reg_activation27_18_1), .reg_activation22(reg_activation27_18_2), .weight_en(weight_en));
SA22 U27_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_19_1), .partial_sum_in12(reg_psum26_19_2), .weight_in11(reg_weight26_19_1), .weight_in12(reg_weight26_19_2), .activation_in11(reg_activation27_18_1), .activation_in21(reg_activation27_18_2), .reg_partial_sum21(reg_psum27_19_1), .reg_partial_sum22(reg_psum27_19_2), .reg_weight21(reg_weight27_19_1), .reg_weight22(reg_weight27_19_2), .reg_activation12(reg_activation27_19_1), .reg_activation22(reg_activation27_19_2), .weight_en(weight_en));
SA22 U27_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_20_1), .partial_sum_in12(reg_psum26_20_2), .weight_in11(reg_weight26_20_1), .weight_in12(reg_weight26_20_2), .activation_in11(reg_activation27_19_1), .activation_in21(reg_activation27_19_2), .reg_partial_sum21(reg_psum27_20_1), .reg_partial_sum22(reg_psum27_20_2), .reg_weight21(reg_weight27_20_1), .reg_weight22(reg_weight27_20_2), .reg_activation12(reg_activation27_20_1), .reg_activation22(reg_activation27_20_2), .weight_en(weight_en));
SA22 U27_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_21_1), .partial_sum_in12(reg_psum26_21_2), .weight_in11(reg_weight26_21_1), .weight_in12(reg_weight26_21_2), .activation_in11(reg_activation27_20_1), .activation_in21(reg_activation27_20_2), .reg_partial_sum21(reg_psum27_21_1), .reg_partial_sum22(reg_psum27_21_2), .reg_weight21(reg_weight27_21_1), .reg_weight22(reg_weight27_21_2), .reg_activation12(reg_activation27_21_1), .reg_activation22(reg_activation27_21_2), .weight_en(weight_en));
SA22 U27_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_22_1), .partial_sum_in12(reg_psum26_22_2), .weight_in11(reg_weight26_22_1), .weight_in12(reg_weight26_22_2), .activation_in11(reg_activation27_21_1), .activation_in21(reg_activation27_21_2), .reg_partial_sum21(reg_psum27_22_1), .reg_partial_sum22(reg_psum27_22_2), .reg_weight21(reg_weight27_22_1), .reg_weight22(reg_weight27_22_2), .reg_activation12(reg_activation27_22_1), .reg_activation22(reg_activation27_22_2), .weight_en(weight_en));
SA22 U27_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_23_1), .partial_sum_in12(reg_psum26_23_2), .weight_in11(reg_weight26_23_1), .weight_in12(reg_weight26_23_2), .activation_in11(reg_activation27_22_1), .activation_in21(reg_activation27_22_2), .reg_partial_sum21(reg_psum27_23_1), .reg_partial_sum22(reg_psum27_23_2), .reg_weight21(reg_weight27_23_1), .reg_weight22(reg_weight27_23_2), .reg_activation12(reg_activation27_23_1), .reg_activation22(reg_activation27_23_2), .weight_en(weight_en));
SA22 U27_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_24_1), .partial_sum_in12(reg_psum26_24_2), .weight_in11(reg_weight26_24_1), .weight_in12(reg_weight26_24_2), .activation_in11(reg_activation27_23_1), .activation_in21(reg_activation27_23_2), .reg_partial_sum21(reg_psum27_24_1), .reg_partial_sum22(reg_psum27_24_2), .reg_weight21(reg_weight27_24_1), .reg_weight22(reg_weight27_24_2), .reg_activation12(reg_activation27_24_1), .reg_activation22(reg_activation27_24_2), .weight_en(weight_en));
SA22 U27_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_25_1), .partial_sum_in12(reg_psum26_25_2), .weight_in11(reg_weight26_25_1), .weight_in12(reg_weight26_25_2), .activation_in11(reg_activation27_24_1), .activation_in21(reg_activation27_24_2), .reg_partial_sum21(reg_psum27_25_1), .reg_partial_sum22(reg_psum27_25_2), .reg_weight21(reg_weight27_25_1), .reg_weight22(reg_weight27_25_2), .reg_activation12(reg_activation27_25_1), .reg_activation22(reg_activation27_25_2), .weight_en(weight_en));
SA22 U27_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_26_1), .partial_sum_in12(reg_psum26_26_2), .weight_in11(reg_weight26_26_1), .weight_in12(reg_weight26_26_2), .activation_in11(reg_activation27_25_1), .activation_in21(reg_activation27_25_2), .reg_partial_sum21(reg_psum27_26_1), .reg_partial_sum22(reg_psum27_26_2), .reg_weight21(reg_weight27_26_1), .reg_weight22(reg_weight27_26_2), .reg_activation12(reg_activation27_26_1), .reg_activation22(reg_activation27_26_2), .weight_en(weight_en));
SA22 U27_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_27_1), .partial_sum_in12(reg_psum26_27_2), .weight_in11(reg_weight26_27_1), .weight_in12(reg_weight26_27_2), .activation_in11(reg_activation27_26_1), .activation_in21(reg_activation27_26_2), .reg_partial_sum21(reg_psum27_27_1), .reg_partial_sum22(reg_psum27_27_2), .reg_weight21(reg_weight27_27_1), .reg_weight22(reg_weight27_27_2), .reg_activation12(reg_activation27_27_1), .reg_activation22(reg_activation27_27_2), .weight_en(weight_en));
SA22 U27_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_28_1), .partial_sum_in12(reg_psum26_28_2), .weight_in11(reg_weight26_28_1), .weight_in12(reg_weight26_28_2), .activation_in11(reg_activation27_27_1), .activation_in21(reg_activation27_27_2), .reg_partial_sum21(reg_psum27_28_1), .reg_partial_sum22(reg_psum27_28_2), .reg_weight21(reg_weight27_28_1), .reg_weight22(reg_weight27_28_2), .reg_activation12(reg_activation27_28_1), .reg_activation22(reg_activation27_28_2), .weight_en(weight_en));
SA22 U27_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_29_1), .partial_sum_in12(reg_psum26_29_2), .weight_in11(reg_weight26_29_1), .weight_in12(reg_weight26_29_2), .activation_in11(reg_activation27_28_1), .activation_in21(reg_activation27_28_2), .reg_partial_sum21(reg_psum27_29_1), .reg_partial_sum22(reg_psum27_29_2), .reg_weight21(reg_weight27_29_1), .reg_weight22(reg_weight27_29_2), .reg_activation12(reg_activation27_29_1), .reg_activation22(reg_activation27_29_2), .weight_en(weight_en));
SA22 U27_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_30_1), .partial_sum_in12(reg_psum26_30_2), .weight_in11(reg_weight26_30_1), .weight_in12(reg_weight26_30_2), .activation_in11(reg_activation27_29_1), .activation_in21(reg_activation27_29_2), .reg_partial_sum21(reg_psum27_30_1), .reg_partial_sum22(reg_psum27_30_2), .reg_weight21(reg_weight27_30_1), .reg_weight22(reg_weight27_30_2), .reg_activation12(reg_activation27_30_1), .reg_activation22(reg_activation27_30_2), .weight_en(weight_en));
SA22 U27_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_31_1), .partial_sum_in12(reg_psum26_31_2), .weight_in11(reg_weight26_31_1), .weight_in12(reg_weight26_31_2), .activation_in11(reg_activation27_30_1), .activation_in21(reg_activation27_30_2), .reg_partial_sum21(reg_psum27_31_1), .reg_partial_sum22(reg_psum27_31_2), .reg_weight21(reg_weight27_31_1), .reg_weight22(reg_weight27_31_2), .reg_activation12(reg_activation27_31_1), .reg_activation22(reg_activation27_31_2), .weight_en(weight_en));
SA22 U27_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum26_32_1), .partial_sum_in12(reg_psum26_32_2), .weight_in11(reg_weight26_32_1), .weight_in12(reg_weight26_32_2), .activation_in11(reg_activation27_31_1), .activation_in21(reg_activation27_31_2), .reg_partial_sum21(reg_psum27_32_1), .reg_partial_sum22(reg_psum27_32_2), .reg_weight21(reg_weight27_32_1), .reg_weight22(reg_weight27_32_2), .weight_en(weight_en));
SA22 U28_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_1_1), .partial_sum_in12(reg_psum27_1_2), .weight_in11(reg_weight27_1_1), .weight_in12(reg_weight27_1_2), .activation_in11(in_activation28_1_1), .activation_in21(in_activation28_1_2), .reg_partial_sum21(reg_psum28_1_1), .reg_partial_sum22(reg_psum28_1_2), .reg_weight21(reg_weight28_1_1), .reg_weight22(reg_weight28_1_2), .reg_activation12(reg_activation28_1_1), .reg_activation22(reg_activation28_1_2), .weight_en(weight_en));
SA22 U28_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_2_1), .partial_sum_in12(reg_psum27_2_2), .weight_in11(reg_weight27_2_1), .weight_in12(reg_weight27_2_2), .activation_in11(reg_activation28_1_1), .activation_in21(reg_activation28_1_2), .reg_partial_sum21(reg_psum28_2_1), .reg_partial_sum22(reg_psum28_2_2), .reg_weight21(reg_weight28_2_1), .reg_weight22(reg_weight28_2_2), .reg_activation12(reg_activation28_2_1), .reg_activation22(reg_activation28_2_2), .weight_en(weight_en));
SA22 U28_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_3_1), .partial_sum_in12(reg_psum27_3_2), .weight_in11(reg_weight27_3_1), .weight_in12(reg_weight27_3_2), .activation_in11(reg_activation28_2_1), .activation_in21(reg_activation28_2_2), .reg_partial_sum21(reg_psum28_3_1), .reg_partial_sum22(reg_psum28_3_2), .reg_weight21(reg_weight28_3_1), .reg_weight22(reg_weight28_3_2), .reg_activation12(reg_activation28_3_1), .reg_activation22(reg_activation28_3_2), .weight_en(weight_en));
SA22 U28_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_4_1), .partial_sum_in12(reg_psum27_4_2), .weight_in11(reg_weight27_4_1), .weight_in12(reg_weight27_4_2), .activation_in11(reg_activation28_3_1), .activation_in21(reg_activation28_3_2), .reg_partial_sum21(reg_psum28_4_1), .reg_partial_sum22(reg_psum28_4_2), .reg_weight21(reg_weight28_4_1), .reg_weight22(reg_weight28_4_2), .reg_activation12(reg_activation28_4_1), .reg_activation22(reg_activation28_4_2), .weight_en(weight_en));
SA22 U28_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_5_1), .partial_sum_in12(reg_psum27_5_2), .weight_in11(reg_weight27_5_1), .weight_in12(reg_weight27_5_2), .activation_in11(reg_activation28_4_1), .activation_in21(reg_activation28_4_2), .reg_partial_sum21(reg_psum28_5_1), .reg_partial_sum22(reg_psum28_5_2), .reg_weight21(reg_weight28_5_1), .reg_weight22(reg_weight28_5_2), .reg_activation12(reg_activation28_5_1), .reg_activation22(reg_activation28_5_2), .weight_en(weight_en));
SA22 U28_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_6_1), .partial_sum_in12(reg_psum27_6_2), .weight_in11(reg_weight27_6_1), .weight_in12(reg_weight27_6_2), .activation_in11(reg_activation28_5_1), .activation_in21(reg_activation28_5_2), .reg_partial_sum21(reg_psum28_6_1), .reg_partial_sum22(reg_psum28_6_2), .reg_weight21(reg_weight28_6_1), .reg_weight22(reg_weight28_6_2), .reg_activation12(reg_activation28_6_1), .reg_activation22(reg_activation28_6_2), .weight_en(weight_en));
SA22 U28_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_7_1), .partial_sum_in12(reg_psum27_7_2), .weight_in11(reg_weight27_7_1), .weight_in12(reg_weight27_7_2), .activation_in11(reg_activation28_6_1), .activation_in21(reg_activation28_6_2), .reg_partial_sum21(reg_psum28_7_1), .reg_partial_sum22(reg_psum28_7_2), .reg_weight21(reg_weight28_7_1), .reg_weight22(reg_weight28_7_2), .reg_activation12(reg_activation28_7_1), .reg_activation22(reg_activation28_7_2), .weight_en(weight_en));
SA22 U28_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_8_1), .partial_sum_in12(reg_psum27_8_2), .weight_in11(reg_weight27_8_1), .weight_in12(reg_weight27_8_2), .activation_in11(reg_activation28_7_1), .activation_in21(reg_activation28_7_2), .reg_partial_sum21(reg_psum28_8_1), .reg_partial_sum22(reg_psum28_8_2), .reg_weight21(reg_weight28_8_1), .reg_weight22(reg_weight28_8_2), .reg_activation12(reg_activation28_8_1), .reg_activation22(reg_activation28_8_2), .weight_en(weight_en));
SA22 U28_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_9_1), .partial_sum_in12(reg_psum27_9_2), .weight_in11(reg_weight27_9_1), .weight_in12(reg_weight27_9_2), .activation_in11(reg_activation28_8_1), .activation_in21(reg_activation28_8_2), .reg_partial_sum21(reg_psum28_9_1), .reg_partial_sum22(reg_psum28_9_2), .reg_weight21(reg_weight28_9_1), .reg_weight22(reg_weight28_9_2), .reg_activation12(reg_activation28_9_1), .reg_activation22(reg_activation28_9_2), .weight_en(weight_en));
SA22 U28_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_10_1), .partial_sum_in12(reg_psum27_10_2), .weight_in11(reg_weight27_10_1), .weight_in12(reg_weight27_10_2), .activation_in11(reg_activation28_9_1), .activation_in21(reg_activation28_9_2), .reg_partial_sum21(reg_psum28_10_1), .reg_partial_sum22(reg_psum28_10_2), .reg_weight21(reg_weight28_10_1), .reg_weight22(reg_weight28_10_2), .reg_activation12(reg_activation28_10_1), .reg_activation22(reg_activation28_10_2), .weight_en(weight_en));
SA22 U28_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_11_1), .partial_sum_in12(reg_psum27_11_2), .weight_in11(reg_weight27_11_1), .weight_in12(reg_weight27_11_2), .activation_in11(reg_activation28_10_1), .activation_in21(reg_activation28_10_2), .reg_partial_sum21(reg_psum28_11_1), .reg_partial_sum22(reg_psum28_11_2), .reg_weight21(reg_weight28_11_1), .reg_weight22(reg_weight28_11_2), .reg_activation12(reg_activation28_11_1), .reg_activation22(reg_activation28_11_2), .weight_en(weight_en));
SA22 U28_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_12_1), .partial_sum_in12(reg_psum27_12_2), .weight_in11(reg_weight27_12_1), .weight_in12(reg_weight27_12_2), .activation_in11(reg_activation28_11_1), .activation_in21(reg_activation28_11_2), .reg_partial_sum21(reg_psum28_12_1), .reg_partial_sum22(reg_psum28_12_2), .reg_weight21(reg_weight28_12_1), .reg_weight22(reg_weight28_12_2), .reg_activation12(reg_activation28_12_1), .reg_activation22(reg_activation28_12_2), .weight_en(weight_en));
SA22 U28_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_13_1), .partial_sum_in12(reg_psum27_13_2), .weight_in11(reg_weight27_13_1), .weight_in12(reg_weight27_13_2), .activation_in11(reg_activation28_12_1), .activation_in21(reg_activation28_12_2), .reg_partial_sum21(reg_psum28_13_1), .reg_partial_sum22(reg_psum28_13_2), .reg_weight21(reg_weight28_13_1), .reg_weight22(reg_weight28_13_2), .reg_activation12(reg_activation28_13_1), .reg_activation22(reg_activation28_13_2), .weight_en(weight_en));
SA22 U28_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_14_1), .partial_sum_in12(reg_psum27_14_2), .weight_in11(reg_weight27_14_1), .weight_in12(reg_weight27_14_2), .activation_in11(reg_activation28_13_1), .activation_in21(reg_activation28_13_2), .reg_partial_sum21(reg_psum28_14_1), .reg_partial_sum22(reg_psum28_14_2), .reg_weight21(reg_weight28_14_1), .reg_weight22(reg_weight28_14_2), .reg_activation12(reg_activation28_14_1), .reg_activation22(reg_activation28_14_2), .weight_en(weight_en));
SA22 U28_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_15_1), .partial_sum_in12(reg_psum27_15_2), .weight_in11(reg_weight27_15_1), .weight_in12(reg_weight27_15_2), .activation_in11(reg_activation28_14_1), .activation_in21(reg_activation28_14_2), .reg_partial_sum21(reg_psum28_15_1), .reg_partial_sum22(reg_psum28_15_2), .reg_weight21(reg_weight28_15_1), .reg_weight22(reg_weight28_15_2), .reg_activation12(reg_activation28_15_1), .reg_activation22(reg_activation28_15_2), .weight_en(weight_en));
SA22 U28_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_16_1), .partial_sum_in12(reg_psum27_16_2), .weight_in11(reg_weight27_16_1), .weight_in12(reg_weight27_16_2), .activation_in11(reg_activation28_15_1), .activation_in21(reg_activation28_15_2), .reg_partial_sum21(reg_psum28_16_1), .reg_partial_sum22(reg_psum28_16_2), .reg_weight21(reg_weight28_16_1), .reg_weight22(reg_weight28_16_2), .reg_activation12(reg_activation28_16_1), .reg_activation22(reg_activation28_16_2), .weight_en(weight_en));
SA22 U28_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_17_1), .partial_sum_in12(reg_psum27_17_2), .weight_in11(reg_weight27_17_1), .weight_in12(reg_weight27_17_2), .activation_in11(reg_activation28_16_1), .activation_in21(reg_activation28_16_2), .reg_partial_sum21(reg_psum28_17_1), .reg_partial_sum22(reg_psum28_17_2), .reg_weight21(reg_weight28_17_1), .reg_weight22(reg_weight28_17_2), .reg_activation12(reg_activation28_17_1), .reg_activation22(reg_activation28_17_2), .weight_en(weight_en));
SA22 U28_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_18_1), .partial_sum_in12(reg_psum27_18_2), .weight_in11(reg_weight27_18_1), .weight_in12(reg_weight27_18_2), .activation_in11(reg_activation28_17_1), .activation_in21(reg_activation28_17_2), .reg_partial_sum21(reg_psum28_18_1), .reg_partial_sum22(reg_psum28_18_2), .reg_weight21(reg_weight28_18_1), .reg_weight22(reg_weight28_18_2), .reg_activation12(reg_activation28_18_1), .reg_activation22(reg_activation28_18_2), .weight_en(weight_en));
SA22 U28_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_19_1), .partial_sum_in12(reg_psum27_19_2), .weight_in11(reg_weight27_19_1), .weight_in12(reg_weight27_19_2), .activation_in11(reg_activation28_18_1), .activation_in21(reg_activation28_18_2), .reg_partial_sum21(reg_psum28_19_1), .reg_partial_sum22(reg_psum28_19_2), .reg_weight21(reg_weight28_19_1), .reg_weight22(reg_weight28_19_2), .reg_activation12(reg_activation28_19_1), .reg_activation22(reg_activation28_19_2), .weight_en(weight_en));
SA22 U28_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_20_1), .partial_sum_in12(reg_psum27_20_2), .weight_in11(reg_weight27_20_1), .weight_in12(reg_weight27_20_2), .activation_in11(reg_activation28_19_1), .activation_in21(reg_activation28_19_2), .reg_partial_sum21(reg_psum28_20_1), .reg_partial_sum22(reg_psum28_20_2), .reg_weight21(reg_weight28_20_1), .reg_weight22(reg_weight28_20_2), .reg_activation12(reg_activation28_20_1), .reg_activation22(reg_activation28_20_2), .weight_en(weight_en));
SA22 U28_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_21_1), .partial_sum_in12(reg_psum27_21_2), .weight_in11(reg_weight27_21_1), .weight_in12(reg_weight27_21_2), .activation_in11(reg_activation28_20_1), .activation_in21(reg_activation28_20_2), .reg_partial_sum21(reg_psum28_21_1), .reg_partial_sum22(reg_psum28_21_2), .reg_weight21(reg_weight28_21_1), .reg_weight22(reg_weight28_21_2), .reg_activation12(reg_activation28_21_1), .reg_activation22(reg_activation28_21_2), .weight_en(weight_en));
SA22 U28_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_22_1), .partial_sum_in12(reg_psum27_22_2), .weight_in11(reg_weight27_22_1), .weight_in12(reg_weight27_22_2), .activation_in11(reg_activation28_21_1), .activation_in21(reg_activation28_21_2), .reg_partial_sum21(reg_psum28_22_1), .reg_partial_sum22(reg_psum28_22_2), .reg_weight21(reg_weight28_22_1), .reg_weight22(reg_weight28_22_2), .reg_activation12(reg_activation28_22_1), .reg_activation22(reg_activation28_22_2), .weight_en(weight_en));
SA22 U28_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_23_1), .partial_sum_in12(reg_psum27_23_2), .weight_in11(reg_weight27_23_1), .weight_in12(reg_weight27_23_2), .activation_in11(reg_activation28_22_1), .activation_in21(reg_activation28_22_2), .reg_partial_sum21(reg_psum28_23_1), .reg_partial_sum22(reg_psum28_23_2), .reg_weight21(reg_weight28_23_1), .reg_weight22(reg_weight28_23_2), .reg_activation12(reg_activation28_23_1), .reg_activation22(reg_activation28_23_2), .weight_en(weight_en));
SA22 U28_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_24_1), .partial_sum_in12(reg_psum27_24_2), .weight_in11(reg_weight27_24_1), .weight_in12(reg_weight27_24_2), .activation_in11(reg_activation28_23_1), .activation_in21(reg_activation28_23_2), .reg_partial_sum21(reg_psum28_24_1), .reg_partial_sum22(reg_psum28_24_2), .reg_weight21(reg_weight28_24_1), .reg_weight22(reg_weight28_24_2), .reg_activation12(reg_activation28_24_1), .reg_activation22(reg_activation28_24_2), .weight_en(weight_en));
SA22 U28_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_25_1), .partial_sum_in12(reg_psum27_25_2), .weight_in11(reg_weight27_25_1), .weight_in12(reg_weight27_25_2), .activation_in11(reg_activation28_24_1), .activation_in21(reg_activation28_24_2), .reg_partial_sum21(reg_psum28_25_1), .reg_partial_sum22(reg_psum28_25_2), .reg_weight21(reg_weight28_25_1), .reg_weight22(reg_weight28_25_2), .reg_activation12(reg_activation28_25_1), .reg_activation22(reg_activation28_25_2), .weight_en(weight_en));
SA22 U28_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_26_1), .partial_sum_in12(reg_psum27_26_2), .weight_in11(reg_weight27_26_1), .weight_in12(reg_weight27_26_2), .activation_in11(reg_activation28_25_1), .activation_in21(reg_activation28_25_2), .reg_partial_sum21(reg_psum28_26_1), .reg_partial_sum22(reg_psum28_26_2), .reg_weight21(reg_weight28_26_1), .reg_weight22(reg_weight28_26_2), .reg_activation12(reg_activation28_26_1), .reg_activation22(reg_activation28_26_2), .weight_en(weight_en));
SA22 U28_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_27_1), .partial_sum_in12(reg_psum27_27_2), .weight_in11(reg_weight27_27_1), .weight_in12(reg_weight27_27_2), .activation_in11(reg_activation28_26_1), .activation_in21(reg_activation28_26_2), .reg_partial_sum21(reg_psum28_27_1), .reg_partial_sum22(reg_psum28_27_2), .reg_weight21(reg_weight28_27_1), .reg_weight22(reg_weight28_27_2), .reg_activation12(reg_activation28_27_1), .reg_activation22(reg_activation28_27_2), .weight_en(weight_en));
SA22 U28_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_28_1), .partial_sum_in12(reg_psum27_28_2), .weight_in11(reg_weight27_28_1), .weight_in12(reg_weight27_28_2), .activation_in11(reg_activation28_27_1), .activation_in21(reg_activation28_27_2), .reg_partial_sum21(reg_psum28_28_1), .reg_partial_sum22(reg_psum28_28_2), .reg_weight21(reg_weight28_28_1), .reg_weight22(reg_weight28_28_2), .reg_activation12(reg_activation28_28_1), .reg_activation22(reg_activation28_28_2), .weight_en(weight_en));
SA22 U28_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_29_1), .partial_sum_in12(reg_psum27_29_2), .weight_in11(reg_weight27_29_1), .weight_in12(reg_weight27_29_2), .activation_in11(reg_activation28_28_1), .activation_in21(reg_activation28_28_2), .reg_partial_sum21(reg_psum28_29_1), .reg_partial_sum22(reg_psum28_29_2), .reg_weight21(reg_weight28_29_1), .reg_weight22(reg_weight28_29_2), .reg_activation12(reg_activation28_29_1), .reg_activation22(reg_activation28_29_2), .weight_en(weight_en));
SA22 U28_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_30_1), .partial_sum_in12(reg_psum27_30_2), .weight_in11(reg_weight27_30_1), .weight_in12(reg_weight27_30_2), .activation_in11(reg_activation28_29_1), .activation_in21(reg_activation28_29_2), .reg_partial_sum21(reg_psum28_30_1), .reg_partial_sum22(reg_psum28_30_2), .reg_weight21(reg_weight28_30_1), .reg_weight22(reg_weight28_30_2), .reg_activation12(reg_activation28_30_1), .reg_activation22(reg_activation28_30_2), .weight_en(weight_en));
SA22 U28_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_31_1), .partial_sum_in12(reg_psum27_31_2), .weight_in11(reg_weight27_31_1), .weight_in12(reg_weight27_31_2), .activation_in11(reg_activation28_30_1), .activation_in21(reg_activation28_30_2), .reg_partial_sum21(reg_psum28_31_1), .reg_partial_sum22(reg_psum28_31_2), .reg_weight21(reg_weight28_31_1), .reg_weight22(reg_weight28_31_2), .reg_activation12(reg_activation28_31_1), .reg_activation22(reg_activation28_31_2), .weight_en(weight_en));
SA22 U28_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum27_32_1), .partial_sum_in12(reg_psum27_32_2), .weight_in11(reg_weight27_32_1), .weight_in12(reg_weight27_32_2), .activation_in11(reg_activation28_31_1), .activation_in21(reg_activation28_31_2), .reg_partial_sum21(reg_psum28_32_1), .reg_partial_sum22(reg_psum28_32_2), .reg_weight21(reg_weight28_32_1), .reg_weight22(reg_weight28_32_2), .weight_en(weight_en));
SA22 U29_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_1_1), .partial_sum_in12(reg_psum28_1_2), .weight_in11(reg_weight28_1_1), .weight_in12(reg_weight28_1_2), .activation_in11(in_activation29_1_1), .activation_in21(in_activation29_1_2), .reg_partial_sum21(reg_psum29_1_1), .reg_partial_sum22(reg_psum29_1_2), .reg_weight21(reg_weight29_1_1), .reg_weight22(reg_weight29_1_2), .reg_activation12(reg_activation29_1_1), .reg_activation22(reg_activation29_1_2), .weight_en(weight_en));
SA22 U29_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_2_1), .partial_sum_in12(reg_psum28_2_2), .weight_in11(reg_weight28_2_1), .weight_in12(reg_weight28_2_2), .activation_in11(reg_activation29_1_1), .activation_in21(reg_activation29_1_2), .reg_partial_sum21(reg_psum29_2_1), .reg_partial_sum22(reg_psum29_2_2), .reg_weight21(reg_weight29_2_1), .reg_weight22(reg_weight29_2_2), .reg_activation12(reg_activation29_2_1), .reg_activation22(reg_activation29_2_2), .weight_en(weight_en));
SA22 U29_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_3_1), .partial_sum_in12(reg_psum28_3_2), .weight_in11(reg_weight28_3_1), .weight_in12(reg_weight28_3_2), .activation_in11(reg_activation29_2_1), .activation_in21(reg_activation29_2_2), .reg_partial_sum21(reg_psum29_3_1), .reg_partial_sum22(reg_psum29_3_2), .reg_weight21(reg_weight29_3_1), .reg_weight22(reg_weight29_3_2), .reg_activation12(reg_activation29_3_1), .reg_activation22(reg_activation29_3_2), .weight_en(weight_en));
SA22 U29_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_4_1), .partial_sum_in12(reg_psum28_4_2), .weight_in11(reg_weight28_4_1), .weight_in12(reg_weight28_4_2), .activation_in11(reg_activation29_3_1), .activation_in21(reg_activation29_3_2), .reg_partial_sum21(reg_psum29_4_1), .reg_partial_sum22(reg_psum29_4_2), .reg_weight21(reg_weight29_4_1), .reg_weight22(reg_weight29_4_2), .reg_activation12(reg_activation29_4_1), .reg_activation22(reg_activation29_4_2), .weight_en(weight_en));
SA22 U29_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_5_1), .partial_sum_in12(reg_psum28_5_2), .weight_in11(reg_weight28_5_1), .weight_in12(reg_weight28_5_2), .activation_in11(reg_activation29_4_1), .activation_in21(reg_activation29_4_2), .reg_partial_sum21(reg_psum29_5_1), .reg_partial_sum22(reg_psum29_5_2), .reg_weight21(reg_weight29_5_1), .reg_weight22(reg_weight29_5_2), .reg_activation12(reg_activation29_5_1), .reg_activation22(reg_activation29_5_2), .weight_en(weight_en));
SA22 U29_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_6_1), .partial_sum_in12(reg_psum28_6_2), .weight_in11(reg_weight28_6_1), .weight_in12(reg_weight28_6_2), .activation_in11(reg_activation29_5_1), .activation_in21(reg_activation29_5_2), .reg_partial_sum21(reg_psum29_6_1), .reg_partial_sum22(reg_psum29_6_2), .reg_weight21(reg_weight29_6_1), .reg_weight22(reg_weight29_6_2), .reg_activation12(reg_activation29_6_1), .reg_activation22(reg_activation29_6_2), .weight_en(weight_en));
SA22 U29_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_7_1), .partial_sum_in12(reg_psum28_7_2), .weight_in11(reg_weight28_7_1), .weight_in12(reg_weight28_7_2), .activation_in11(reg_activation29_6_1), .activation_in21(reg_activation29_6_2), .reg_partial_sum21(reg_psum29_7_1), .reg_partial_sum22(reg_psum29_7_2), .reg_weight21(reg_weight29_7_1), .reg_weight22(reg_weight29_7_2), .reg_activation12(reg_activation29_7_1), .reg_activation22(reg_activation29_7_2), .weight_en(weight_en));
SA22 U29_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_8_1), .partial_sum_in12(reg_psum28_8_2), .weight_in11(reg_weight28_8_1), .weight_in12(reg_weight28_8_2), .activation_in11(reg_activation29_7_1), .activation_in21(reg_activation29_7_2), .reg_partial_sum21(reg_psum29_8_1), .reg_partial_sum22(reg_psum29_8_2), .reg_weight21(reg_weight29_8_1), .reg_weight22(reg_weight29_8_2), .reg_activation12(reg_activation29_8_1), .reg_activation22(reg_activation29_8_2), .weight_en(weight_en));
SA22 U29_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_9_1), .partial_sum_in12(reg_psum28_9_2), .weight_in11(reg_weight28_9_1), .weight_in12(reg_weight28_9_2), .activation_in11(reg_activation29_8_1), .activation_in21(reg_activation29_8_2), .reg_partial_sum21(reg_psum29_9_1), .reg_partial_sum22(reg_psum29_9_2), .reg_weight21(reg_weight29_9_1), .reg_weight22(reg_weight29_9_2), .reg_activation12(reg_activation29_9_1), .reg_activation22(reg_activation29_9_2), .weight_en(weight_en));
SA22 U29_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_10_1), .partial_sum_in12(reg_psum28_10_2), .weight_in11(reg_weight28_10_1), .weight_in12(reg_weight28_10_2), .activation_in11(reg_activation29_9_1), .activation_in21(reg_activation29_9_2), .reg_partial_sum21(reg_psum29_10_1), .reg_partial_sum22(reg_psum29_10_2), .reg_weight21(reg_weight29_10_1), .reg_weight22(reg_weight29_10_2), .reg_activation12(reg_activation29_10_1), .reg_activation22(reg_activation29_10_2), .weight_en(weight_en));
SA22 U29_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_11_1), .partial_sum_in12(reg_psum28_11_2), .weight_in11(reg_weight28_11_1), .weight_in12(reg_weight28_11_2), .activation_in11(reg_activation29_10_1), .activation_in21(reg_activation29_10_2), .reg_partial_sum21(reg_psum29_11_1), .reg_partial_sum22(reg_psum29_11_2), .reg_weight21(reg_weight29_11_1), .reg_weight22(reg_weight29_11_2), .reg_activation12(reg_activation29_11_1), .reg_activation22(reg_activation29_11_2), .weight_en(weight_en));
SA22 U29_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_12_1), .partial_sum_in12(reg_psum28_12_2), .weight_in11(reg_weight28_12_1), .weight_in12(reg_weight28_12_2), .activation_in11(reg_activation29_11_1), .activation_in21(reg_activation29_11_2), .reg_partial_sum21(reg_psum29_12_1), .reg_partial_sum22(reg_psum29_12_2), .reg_weight21(reg_weight29_12_1), .reg_weight22(reg_weight29_12_2), .reg_activation12(reg_activation29_12_1), .reg_activation22(reg_activation29_12_2), .weight_en(weight_en));
SA22 U29_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_13_1), .partial_sum_in12(reg_psum28_13_2), .weight_in11(reg_weight28_13_1), .weight_in12(reg_weight28_13_2), .activation_in11(reg_activation29_12_1), .activation_in21(reg_activation29_12_2), .reg_partial_sum21(reg_psum29_13_1), .reg_partial_sum22(reg_psum29_13_2), .reg_weight21(reg_weight29_13_1), .reg_weight22(reg_weight29_13_2), .reg_activation12(reg_activation29_13_1), .reg_activation22(reg_activation29_13_2), .weight_en(weight_en));
SA22 U29_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_14_1), .partial_sum_in12(reg_psum28_14_2), .weight_in11(reg_weight28_14_1), .weight_in12(reg_weight28_14_2), .activation_in11(reg_activation29_13_1), .activation_in21(reg_activation29_13_2), .reg_partial_sum21(reg_psum29_14_1), .reg_partial_sum22(reg_psum29_14_2), .reg_weight21(reg_weight29_14_1), .reg_weight22(reg_weight29_14_2), .reg_activation12(reg_activation29_14_1), .reg_activation22(reg_activation29_14_2), .weight_en(weight_en));
SA22 U29_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_15_1), .partial_sum_in12(reg_psum28_15_2), .weight_in11(reg_weight28_15_1), .weight_in12(reg_weight28_15_2), .activation_in11(reg_activation29_14_1), .activation_in21(reg_activation29_14_2), .reg_partial_sum21(reg_psum29_15_1), .reg_partial_sum22(reg_psum29_15_2), .reg_weight21(reg_weight29_15_1), .reg_weight22(reg_weight29_15_2), .reg_activation12(reg_activation29_15_1), .reg_activation22(reg_activation29_15_2), .weight_en(weight_en));
SA22 U29_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_16_1), .partial_sum_in12(reg_psum28_16_2), .weight_in11(reg_weight28_16_1), .weight_in12(reg_weight28_16_2), .activation_in11(reg_activation29_15_1), .activation_in21(reg_activation29_15_2), .reg_partial_sum21(reg_psum29_16_1), .reg_partial_sum22(reg_psum29_16_2), .reg_weight21(reg_weight29_16_1), .reg_weight22(reg_weight29_16_2), .reg_activation12(reg_activation29_16_1), .reg_activation22(reg_activation29_16_2), .weight_en(weight_en));
SA22 U29_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_17_1), .partial_sum_in12(reg_psum28_17_2), .weight_in11(reg_weight28_17_1), .weight_in12(reg_weight28_17_2), .activation_in11(reg_activation29_16_1), .activation_in21(reg_activation29_16_2), .reg_partial_sum21(reg_psum29_17_1), .reg_partial_sum22(reg_psum29_17_2), .reg_weight21(reg_weight29_17_1), .reg_weight22(reg_weight29_17_2), .reg_activation12(reg_activation29_17_1), .reg_activation22(reg_activation29_17_2), .weight_en(weight_en));
SA22 U29_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_18_1), .partial_sum_in12(reg_psum28_18_2), .weight_in11(reg_weight28_18_1), .weight_in12(reg_weight28_18_2), .activation_in11(reg_activation29_17_1), .activation_in21(reg_activation29_17_2), .reg_partial_sum21(reg_psum29_18_1), .reg_partial_sum22(reg_psum29_18_2), .reg_weight21(reg_weight29_18_1), .reg_weight22(reg_weight29_18_2), .reg_activation12(reg_activation29_18_1), .reg_activation22(reg_activation29_18_2), .weight_en(weight_en));
SA22 U29_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_19_1), .partial_sum_in12(reg_psum28_19_2), .weight_in11(reg_weight28_19_1), .weight_in12(reg_weight28_19_2), .activation_in11(reg_activation29_18_1), .activation_in21(reg_activation29_18_2), .reg_partial_sum21(reg_psum29_19_1), .reg_partial_sum22(reg_psum29_19_2), .reg_weight21(reg_weight29_19_1), .reg_weight22(reg_weight29_19_2), .reg_activation12(reg_activation29_19_1), .reg_activation22(reg_activation29_19_2), .weight_en(weight_en));
SA22 U29_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_20_1), .partial_sum_in12(reg_psum28_20_2), .weight_in11(reg_weight28_20_1), .weight_in12(reg_weight28_20_2), .activation_in11(reg_activation29_19_1), .activation_in21(reg_activation29_19_2), .reg_partial_sum21(reg_psum29_20_1), .reg_partial_sum22(reg_psum29_20_2), .reg_weight21(reg_weight29_20_1), .reg_weight22(reg_weight29_20_2), .reg_activation12(reg_activation29_20_1), .reg_activation22(reg_activation29_20_2), .weight_en(weight_en));
SA22 U29_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_21_1), .partial_sum_in12(reg_psum28_21_2), .weight_in11(reg_weight28_21_1), .weight_in12(reg_weight28_21_2), .activation_in11(reg_activation29_20_1), .activation_in21(reg_activation29_20_2), .reg_partial_sum21(reg_psum29_21_1), .reg_partial_sum22(reg_psum29_21_2), .reg_weight21(reg_weight29_21_1), .reg_weight22(reg_weight29_21_2), .reg_activation12(reg_activation29_21_1), .reg_activation22(reg_activation29_21_2), .weight_en(weight_en));
SA22 U29_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_22_1), .partial_sum_in12(reg_psum28_22_2), .weight_in11(reg_weight28_22_1), .weight_in12(reg_weight28_22_2), .activation_in11(reg_activation29_21_1), .activation_in21(reg_activation29_21_2), .reg_partial_sum21(reg_psum29_22_1), .reg_partial_sum22(reg_psum29_22_2), .reg_weight21(reg_weight29_22_1), .reg_weight22(reg_weight29_22_2), .reg_activation12(reg_activation29_22_1), .reg_activation22(reg_activation29_22_2), .weight_en(weight_en));
SA22 U29_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_23_1), .partial_sum_in12(reg_psum28_23_2), .weight_in11(reg_weight28_23_1), .weight_in12(reg_weight28_23_2), .activation_in11(reg_activation29_22_1), .activation_in21(reg_activation29_22_2), .reg_partial_sum21(reg_psum29_23_1), .reg_partial_sum22(reg_psum29_23_2), .reg_weight21(reg_weight29_23_1), .reg_weight22(reg_weight29_23_2), .reg_activation12(reg_activation29_23_1), .reg_activation22(reg_activation29_23_2), .weight_en(weight_en));
SA22 U29_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_24_1), .partial_sum_in12(reg_psum28_24_2), .weight_in11(reg_weight28_24_1), .weight_in12(reg_weight28_24_2), .activation_in11(reg_activation29_23_1), .activation_in21(reg_activation29_23_2), .reg_partial_sum21(reg_psum29_24_1), .reg_partial_sum22(reg_psum29_24_2), .reg_weight21(reg_weight29_24_1), .reg_weight22(reg_weight29_24_2), .reg_activation12(reg_activation29_24_1), .reg_activation22(reg_activation29_24_2), .weight_en(weight_en));
SA22 U29_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_25_1), .partial_sum_in12(reg_psum28_25_2), .weight_in11(reg_weight28_25_1), .weight_in12(reg_weight28_25_2), .activation_in11(reg_activation29_24_1), .activation_in21(reg_activation29_24_2), .reg_partial_sum21(reg_psum29_25_1), .reg_partial_sum22(reg_psum29_25_2), .reg_weight21(reg_weight29_25_1), .reg_weight22(reg_weight29_25_2), .reg_activation12(reg_activation29_25_1), .reg_activation22(reg_activation29_25_2), .weight_en(weight_en));
SA22 U29_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_26_1), .partial_sum_in12(reg_psum28_26_2), .weight_in11(reg_weight28_26_1), .weight_in12(reg_weight28_26_2), .activation_in11(reg_activation29_25_1), .activation_in21(reg_activation29_25_2), .reg_partial_sum21(reg_psum29_26_1), .reg_partial_sum22(reg_psum29_26_2), .reg_weight21(reg_weight29_26_1), .reg_weight22(reg_weight29_26_2), .reg_activation12(reg_activation29_26_1), .reg_activation22(reg_activation29_26_2), .weight_en(weight_en));
SA22 U29_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_27_1), .partial_sum_in12(reg_psum28_27_2), .weight_in11(reg_weight28_27_1), .weight_in12(reg_weight28_27_2), .activation_in11(reg_activation29_26_1), .activation_in21(reg_activation29_26_2), .reg_partial_sum21(reg_psum29_27_1), .reg_partial_sum22(reg_psum29_27_2), .reg_weight21(reg_weight29_27_1), .reg_weight22(reg_weight29_27_2), .reg_activation12(reg_activation29_27_1), .reg_activation22(reg_activation29_27_2), .weight_en(weight_en));
SA22 U29_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_28_1), .partial_sum_in12(reg_psum28_28_2), .weight_in11(reg_weight28_28_1), .weight_in12(reg_weight28_28_2), .activation_in11(reg_activation29_27_1), .activation_in21(reg_activation29_27_2), .reg_partial_sum21(reg_psum29_28_1), .reg_partial_sum22(reg_psum29_28_2), .reg_weight21(reg_weight29_28_1), .reg_weight22(reg_weight29_28_2), .reg_activation12(reg_activation29_28_1), .reg_activation22(reg_activation29_28_2), .weight_en(weight_en));
SA22 U29_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_29_1), .partial_sum_in12(reg_psum28_29_2), .weight_in11(reg_weight28_29_1), .weight_in12(reg_weight28_29_2), .activation_in11(reg_activation29_28_1), .activation_in21(reg_activation29_28_2), .reg_partial_sum21(reg_psum29_29_1), .reg_partial_sum22(reg_psum29_29_2), .reg_weight21(reg_weight29_29_1), .reg_weight22(reg_weight29_29_2), .reg_activation12(reg_activation29_29_1), .reg_activation22(reg_activation29_29_2), .weight_en(weight_en));
SA22 U29_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_30_1), .partial_sum_in12(reg_psum28_30_2), .weight_in11(reg_weight28_30_1), .weight_in12(reg_weight28_30_2), .activation_in11(reg_activation29_29_1), .activation_in21(reg_activation29_29_2), .reg_partial_sum21(reg_psum29_30_1), .reg_partial_sum22(reg_psum29_30_2), .reg_weight21(reg_weight29_30_1), .reg_weight22(reg_weight29_30_2), .reg_activation12(reg_activation29_30_1), .reg_activation22(reg_activation29_30_2), .weight_en(weight_en));
SA22 U29_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_31_1), .partial_sum_in12(reg_psum28_31_2), .weight_in11(reg_weight28_31_1), .weight_in12(reg_weight28_31_2), .activation_in11(reg_activation29_30_1), .activation_in21(reg_activation29_30_2), .reg_partial_sum21(reg_psum29_31_1), .reg_partial_sum22(reg_psum29_31_2), .reg_weight21(reg_weight29_31_1), .reg_weight22(reg_weight29_31_2), .reg_activation12(reg_activation29_31_1), .reg_activation22(reg_activation29_31_2), .weight_en(weight_en));
SA22 U29_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum28_32_1), .partial_sum_in12(reg_psum28_32_2), .weight_in11(reg_weight28_32_1), .weight_in12(reg_weight28_32_2), .activation_in11(reg_activation29_31_1), .activation_in21(reg_activation29_31_2), .reg_partial_sum21(reg_psum29_32_1), .reg_partial_sum22(reg_psum29_32_2), .reg_weight21(reg_weight29_32_1), .reg_weight22(reg_weight29_32_2), .weight_en(weight_en));
SA22 U30_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_1_1), .partial_sum_in12(reg_psum29_1_2), .weight_in11(reg_weight29_1_1), .weight_in12(reg_weight29_1_2), .activation_in11(in_activation30_1_1), .activation_in21(in_activation30_1_2), .reg_partial_sum21(reg_psum30_1_1), .reg_partial_sum22(reg_psum30_1_2), .reg_weight21(reg_weight30_1_1), .reg_weight22(reg_weight30_1_2), .reg_activation12(reg_activation30_1_1), .reg_activation22(reg_activation30_1_2), .weight_en(weight_en));
SA22 U30_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_2_1), .partial_sum_in12(reg_psum29_2_2), .weight_in11(reg_weight29_2_1), .weight_in12(reg_weight29_2_2), .activation_in11(reg_activation30_1_1), .activation_in21(reg_activation30_1_2), .reg_partial_sum21(reg_psum30_2_1), .reg_partial_sum22(reg_psum30_2_2), .reg_weight21(reg_weight30_2_1), .reg_weight22(reg_weight30_2_2), .reg_activation12(reg_activation30_2_1), .reg_activation22(reg_activation30_2_2), .weight_en(weight_en));
SA22 U30_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_3_1), .partial_sum_in12(reg_psum29_3_2), .weight_in11(reg_weight29_3_1), .weight_in12(reg_weight29_3_2), .activation_in11(reg_activation30_2_1), .activation_in21(reg_activation30_2_2), .reg_partial_sum21(reg_psum30_3_1), .reg_partial_sum22(reg_psum30_3_2), .reg_weight21(reg_weight30_3_1), .reg_weight22(reg_weight30_3_2), .reg_activation12(reg_activation30_3_1), .reg_activation22(reg_activation30_3_2), .weight_en(weight_en));
SA22 U30_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_4_1), .partial_sum_in12(reg_psum29_4_2), .weight_in11(reg_weight29_4_1), .weight_in12(reg_weight29_4_2), .activation_in11(reg_activation30_3_1), .activation_in21(reg_activation30_3_2), .reg_partial_sum21(reg_psum30_4_1), .reg_partial_sum22(reg_psum30_4_2), .reg_weight21(reg_weight30_4_1), .reg_weight22(reg_weight30_4_2), .reg_activation12(reg_activation30_4_1), .reg_activation22(reg_activation30_4_2), .weight_en(weight_en));
SA22 U30_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_5_1), .partial_sum_in12(reg_psum29_5_2), .weight_in11(reg_weight29_5_1), .weight_in12(reg_weight29_5_2), .activation_in11(reg_activation30_4_1), .activation_in21(reg_activation30_4_2), .reg_partial_sum21(reg_psum30_5_1), .reg_partial_sum22(reg_psum30_5_2), .reg_weight21(reg_weight30_5_1), .reg_weight22(reg_weight30_5_2), .reg_activation12(reg_activation30_5_1), .reg_activation22(reg_activation30_5_2), .weight_en(weight_en));
SA22 U30_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_6_1), .partial_sum_in12(reg_psum29_6_2), .weight_in11(reg_weight29_6_1), .weight_in12(reg_weight29_6_2), .activation_in11(reg_activation30_5_1), .activation_in21(reg_activation30_5_2), .reg_partial_sum21(reg_psum30_6_1), .reg_partial_sum22(reg_psum30_6_2), .reg_weight21(reg_weight30_6_1), .reg_weight22(reg_weight30_6_2), .reg_activation12(reg_activation30_6_1), .reg_activation22(reg_activation30_6_2), .weight_en(weight_en));
SA22 U30_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_7_1), .partial_sum_in12(reg_psum29_7_2), .weight_in11(reg_weight29_7_1), .weight_in12(reg_weight29_7_2), .activation_in11(reg_activation30_6_1), .activation_in21(reg_activation30_6_2), .reg_partial_sum21(reg_psum30_7_1), .reg_partial_sum22(reg_psum30_7_2), .reg_weight21(reg_weight30_7_1), .reg_weight22(reg_weight30_7_2), .reg_activation12(reg_activation30_7_1), .reg_activation22(reg_activation30_7_2), .weight_en(weight_en));
SA22 U30_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_8_1), .partial_sum_in12(reg_psum29_8_2), .weight_in11(reg_weight29_8_1), .weight_in12(reg_weight29_8_2), .activation_in11(reg_activation30_7_1), .activation_in21(reg_activation30_7_2), .reg_partial_sum21(reg_psum30_8_1), .reg_partial_sum22(reg_psum30_8_2), .reg_weight21(reg_weight30_8_1), .reg_weight22(reg_weight30_8_2), .reg_activation12(reg_activation30_8_1), .reg_activation22(reg_activation30_8_2), .weight_en(weight_en));
SA22 U30_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_9_1), .partial_sum_in12(reg_psum29_9_2), .weight_in11(reg_weight29_9_1), .weight_in12(reg_weight29_9_2), .activation_in11(reg_activation30_8_1), .activation_in21(reg_activation30_8_2), .reg_partial_sum21(reg_psum30_9_1), .reg_partial_sum22(reg_psum30_9_2), .reg_weight21(reg_weight30_9_1), .reg_weight22(reg_weight30_9_2), .reg_activation12(reg_activation30_9_1), .reg_activation22(reg_activation30_9_2), .weight_en(weight_en));
SA22 U30_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_10_1), .partial_sum_in12(reg_psum29_10_2), .weight_in11(reg_weight29_10_1), .weight_in12(reg_weight29_10_2), .activation_in11(reg_activation30_9_1), .activation_in21(reg_activation30_9_2), .reg_partial_sum21(reg_psum30_10_1), .reg_partial_sum22(reg_psum30_10_2), .reg_weight21(reg_weight30_10_1), .reg_weight22(reg_weight30_10_2), .reg_activation12(reg_activation30_10_1), .reg_activation22(reg_activation30_10_2), .weight_en(weight_en));
SA22 U30_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_11_1), .partial_sum_in12(reg_psum29_11_2), .weight_in11(reg_weight29_11_1), .weight_in12(reg_weight29_11_2), .activation_in11(reg_activation30_10_1), .activation_in21(reg_activation30_10_2), .reg_partial_sum21(reg_psum30_11_1), .reg_partial_sum22(reg_psum30_11_2), .reg_weight21(reg_weight30_11_1), .reg_weight22(reg_weight30_11_2), .reg_activation12(reg_activation30_11_1), .reg_activation22(reg_activation30_11_2), .weight_en(weight_en));
SA22 U30_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_12_1), .partial_sum_in12(reg_psum29_12_2), .weight_in11(reg_weight29_12_1), .weight_in12(reg_weight29_12_2), .activation_in11(reg_activation30_11_1), .activation_in21(reg_activation30_11_2), .reg_partial_sum21(reg_psum30_12_1), .reg_partial_sum22(reg_psum30_12_2), .reg_weight21(reg_weight30_12_1), .reg_weight22(reg_weight30_12_2), .reg_activation12(reg_activation30_12_1), .reg_activation22(reg_activation30_12_2), .weight_en(weight_en));
SA22 U30_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_13_1), .partial_sum_in12(reg_psum29_13_2), .weight_in11(reg_weight29_13_1), .weight_in12(reg_weight29_13_2), .activation_in11(reg_activation30_12_1), .activation_in21(reg_activation30_12_2), .reg_partial_sum21(reg_psum30_13_1), .reg_partial_sum22(reg_psum30_13_2), .reg_weight21(reg_weight30_13_1), .reg_weight22(reg_weight30_13_2), .reg_activation12(reg_activation30_13_1), .reg_activation22(reg_activation30_13_2), .weight_en(weight_en));
SA22 U30_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_14_1), .partial_sum_in12(reg_psum29_14_2), .weight_in11(reg_weight29_14_1), .weight_in12(reg_weight29_14_2), .activation_in11(reg_activation30_13_1), .activation_in21(reg_activation30_13_2), .reg_partial_sum21(reg_psum30_14_1), .reg_partial_sum22(reg_psum30_14_2), .reg_weight21(reg_weight30_14_1), .reg_weight22(reg_weight30_14_2), .reg_activation12(reg_activation30_14_1), .reg_activation22(reg_activation30_14_2), .weight_en(weight_en));
SA22 U30_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_15_1), .partial_sum_in12(reg_psum29_15_2), .weight_in11(reg_weight29_15_1), .weight_in12(reg_weight29_15_2), .activation_in11(reg_activation30_14_1), .activation_in21(reg_activation30_14_2), .reg_partial_sum21(reg_psum30_15_1), .reg_partial_sum22(reg_psum30_15_2), .reg_weight21(reg_weight30_15_1), .reg_weight22(reg_weight30_15_2), .reg_activation12(reg_activation30_15_1), .reg_activation22(reg_activation30_15_2), .weight_en(weight_en));
SA22 U30_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_16_1), .partial_sum_in12(reg_psum29_16_2), .weight_in11(reg_weight29_16_1), .weight_in12(reg_weight29_16_2), .activation_in11(reg_activation30_15_1), .activation_in21(reg_activation30_15_2), .reg_partial_sum21(reg_psum30_16_1), .reg_partial_sum22(reg_psum30_16_2), .reg_weight21(reg_weight30_16_1), .reg_weight22(reg_weight30_16_2), .reg_activation12(reg_activation30_16_1), .reg_activation22(reg_activation30_16_2), .weight_en(weight_en));
SA22 U30_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_17_1), .partial_sum_in12(reg_psum29_17_2), .weight_in11(reg_weight29_17_1), .weight_in12(reg_weight29_17_2), .activation_in11(reg_activation30_16_1), .activation_in21(reg_activation30_16_2), .reg_partial_sum21(reg_psum30_17_1), .reg_partial_sum22(reg_psum30_17_2), .reg_weight21(reg_weight30_17_1), .reg_weight22(reg_weight30_17_2), .reg_activation12(reg_activation30_17_1), .reg_activation22(reg_activation30_17_2), .weight_en(weight_en));
SA22 U30_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_18_1), .partial_sum_in12(reg_psum29_18_2), .weight_in11(reg_weight29_18_1), .weight_in12(reg_weight29_18_2), .activation_in11(reg_activation30_17_1), .activation_in21(reg_activation30_17_2), .reg_partial_sum21(reg_psum30_18_1), .reg_partial_sum22(reg_psum30_18_2), .reg_weight21(reg_weight30_18_1), .reg_weight22(reg_weight30_18_2), .reg_activation12(reg_activation30_18_1), .reg_activation22(reg_activation30_18_2), .weight_en(weight_en));
SA22 U30_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_19_1), .partial_sum_in12(reg_psum29_19_2), .weight_in11(reg_weight29_19_1), .weight_in12(reg_weight29_19_2), .activation_in11(reg_activation30_18_1), .activation_in21(reg_activation30_18_2), .reg_partial_sum21(reg_psum30_19_1), .reg_partial_sum22(reg_psum30_19_2), .reg_weight21(reg_weight30_19_1), .reg_weight22(reg_weight30_19_2), .reg_activation12(reg_activation30_19_1), .reg_activation22(reg_activation30_19_2), .weight_en(weight_en));
SA22 U30_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_20_1), .partial_sum_in12(reg_psum29_20_2), .weight_in11(reg_weight29_20_1), .weight_in12(reg_weight29_20_2), .activation_in11(reg_activation30_19_1), .activation_in21(reg_activation30_19_2), .reg_partial_sum21(reg_psum30_20_1), .reg_partial_sum22(reg_psum30_20_2), .reg_weight21(reg_weight30_20_1), .reg_weight22(reg_weight30_20_2), .reg_activation12(reg_activation30_20_1), .reg_activation22(reg_activation30_20_2), .weight_en(weight_en));
SA22 U30_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_21_1), .partial_sum_in12(reg_psum29_21_2), .weight_in11(reg_weight29_21_1), .weight_in12(reg_weight29_21_2), .activation_in11(reg_activation30_20_1), .activation_in21(reg_activation30_20_2), .reg_partial_sum21(reg_psum30_21_1), .reg_partial_sum22(reg_psum30_21_2), .reg_weight21(reg_weight30_21_1), .reg_weight22(reg_weight30_21_2), .reg_activation12(reg_activation30_21_1), .reg_activation22(reg_activation30_21_2), .weight_en(weight_en));
SA22 U30_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_22_1), .partial_sum_in12(reg_psum29_22_2), .weight_in11(reg_weight29_22_1), .weight_in12(reg_weight29_22_2), .activation_in11(reg_activation30_21_1), .activation_in21(reg_activation30_21_2), .reg_partial_sum21(reg_psum30_22_1), .reg_partial_sum22(reg_psum30_22_2), .reg_weight21(reg_weight30_22_1), .reg_weight22(reg_weight30_22_2), .reg_activation12(reg_activation30_22_1), .reg_activation22(reg_activation30_22_2), .weight_en(weight_en));
SA22 U30_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_23_1), .partial_sum_in12(reg_psum29_23_2), .weight_in11(reg_weight29_23_1), .weight_in12(reg_weight29_23_2), .activation_in11(reg_activation30_22_1), .activation_in21(reg_activation30_22_2), .reg_partial_sum21(reg_psum30_23_1), .reg_partial_sum22(reg_psum30_23_2), .reg_weight21(reg_weight30_23_1), .reg_weight22(reg_weight30_23_2), .reg_activation12(reg_activation30_23_1), .reg_activation22(reg_activation30_23_2), .weight_en(weight_en));
SA22 U30_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_24_1), .partial_sum_in12(reg_psum29_24_2), .weight_in11(reg_weight29_24_1), .weight_in12(reg_weight29_24_2), .activation_in11(reg_activation30_23_1), .activation_in21(reg_activation30_23_2), .reg_partial_sum21(reg_psum30_24_1), .reg_partial_sum22(reg_psum30_24_2), .reg_weight21(reg_weight30_24_1), .reg_weight22(reg_weight30_24_2), .reg_activation12(reg_activation30_24_1), .reg_activation22(reg_activation30_24_2), .weight_en(weight_en));
SA22 U30_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_25_1), .partial_sum_in12(reg_psum29_25_2), .weight_in11(reg_weight29_25_1), .weight_in12(reg_weight29_25_2), .activation_in11(reg_activation30_24_1), .activation_in21(reg_activation30_24_2), .reg_partial_sum21(reg_psum30_25_1), .reg_partial_sum22(reg_psum30_25_2), .reg_weight21(reg_weight30_25_1), .reg_weight22(reg_weight30_25_2), .reg_activation12(reg_activation30_25_1), .reg_activation22(reg_activation30_25_2), .weight_en(weight_en));
SA22 U30_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_26_1), .partial_sum_in12(reg_psum29_26_2), .weight_in11(reg_weight29_26_1), .weight_in12(reg_weight29_26_2), .activation_in11(reg_activation30_25_1), .activation_in21(reg_activation30_25_2), .reg_partial_sum21(reg_psum30_26_1), .reg_partial_sum22(reg_psum30_26_2), .reg_weight21(reg_weight30_26_1), .reg_weight22(reg_weight30_26_2), .reg_activation12(reg_activation30_26_1), .reg_activation22(reg_activation30_26_2), .weight_en(weight_en));
SA22 U30_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_27_1), .partial_sum_in12(reg_psum29_27_2), .weight_in11(reg_weight29_27_1), .weight_in12(reg_weight29_27_2), .activation_in11(reg_activation30_26_1), .activation_in21(reg_activation30_26_2), .reg_partial_sum21(reg_psum30_27_1), .reg_partial_sum22(reg_psum30_27_2), .reg_weight21(reg_weight30_27_1), .reg_weight22(reg_weight30_27_2), .reg_activation12(reg_activation30_27_1), .reg_activation22(reg_activation30_27_2), .weight_en(weight_en));
SA22 U30_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_28_1), .partial_sum_in12(reg_psum29_28_2), .weight_in11(reg_weight29_28_1), .weight_in12(reg_weight29_28_2), .activation_in11(reg_activation30_27_1), .activation_in21(reg_activation30_27_2), .reg_partial_sum21(reg_psum30_28_1), .reg_partial_sum22(reg_psum30_28_2), .reg_weight21(reg_weight30_28_1), .reg_weight22(reg_weight30_28_2), .reg_activation12(reg_activation30_28_1), .reg_activation22(reg_activation30_28_2), .weight_en(weight_en));
SA22 U30_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_29_1), .partial_sum_in12(reg_psum29_29_2), .weight_in11(reg_weight29_29_1), .weight_in12(reg_weight29_29_2), .activation_in11(reg_activation30_28_1), .activation_in21(reg_activation30_28_2), .reg_partial_sum21(reg_psum30_29_1), .reg_partial_sum22(reg_psum30_29_2), .reg_weight21(reg_weight30_29_1), .reg_weight22(reg_weight30_29_2), .reg_activation12(reg_activation30_29_1), .reg_activation22(reg_activation30_29_2), .weight_en(weight_en));
SA22 U30_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_30_1), .partial_sum_in12(reg_psum29_30_2), .weight_in11(reg_weight29_30_1), .weight_in12(reg_weight29_30_2), .activation_in11(reg_activation30_29_1), .activation_in21(reg_activation30_29_2), .reg_partial_sum21(reg_psum30_30_1), .reg_partial_sum22(reg_psum30_30_2), .reg_weight21(reg_weight30_30_1), .reg_weight22(reg_weight30_30_2), .reg_activation12(reg_activation30_30_1), .reg_activation22(reg_activation30_30_2), .weight_en(weight_en));
SA22 U30_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_31_1), .partial_sum_in12(reg_psum29_31_2), .weight_in11(reg_weight29_31_1), .weight_in12(reg_weight29_31_2), .activation_in11(reg_activation30_30_1), .activation_in21(reg_activation30_30_2), .reg_partial_sum21(reg_psum30_31_1), .reg_partial_sum22(reg_psum30_31_2), .reg_weight21(reg_weight30_31_1), .reg_weight22(reg_weight30_31_2), .reg_activation12(reg_activation30_31_1), .reg_activation22(reg_activation30_31_2), .weight_en(weight_en));
SA22 U30_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum29_32_1), .partial_sum_in12(reg_psum29_32_2), .weight_in11(reg_weight29_32_1), .weight_in12(reg_weight29_32_2), .activation_in11(reg_activation30_31_1), .activation_in21(reg_activation30_31_2), .reg_partial_sum21(reg_psum30_32_1), .reg_partial_sum22(reg_psum30_32_2), .reg_weight21(reg_weight30_32_1), .reg_weight22(reg_weight30_32_2), .weight_en(weight_en));
SA22 U31_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_1_1), .partial_sum_in12(reg_psum30_1_2), .weight_in11(reg_weight30_1_1), .weight_in12(reg_weight30_1_2), .activation_in11(in_activation31_1_1), .activation_in21(in_activation31_1_2), .reg_partial_sum21(reg_psum31_1_1), .reg_partial_sum22(reg_psum31_1_2), .reg_weight21(reg_weight31_1_1), .reg_weight22(reg_weight31_1_2), .reg_activation12(reg_activation31_1_1), .reg_activation22(reg_activation31_1_2), .weight_en(weight_en));
SA22 U31_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_2_1), .partial_sum_in12(reg_psum30_2_2), .weight_in11(reg_weight30_2_1), .weight_in12(reg_weight30_2_2), .activation_in11(reg_activation31_1_1), .activation_in21(reg_activation31_1_2), .reg_partial_sum21(reg_psum31_2_1), .reg_partial_sum22(reg_psum31_2_2), .reg_weight21(reg_weight31_2_1), .reg_weight22(reg_weight31_2_2), .reg_activation12(reg_activation31_2_1), .reg_activation22(reg_activation31_2_2), .weight_en(weight_en));
SA22 U31_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_3_1), .partial_sum_in12(reg_psum30_3_2), .weight_in11(reg_weight30_3_1), .weight_in12(reg_weight30_3_2), .activation_in11(reg_activation31_2_1), .activation_in21(reg_activation31_2_2), .reg_partial_sum21(reg_psum31_3_1), .reg_partial_sum22(reg_psum31_3_2), .reg_weight21(reg_weight31_3_1), .reg_weight22(reg_weight31_3_2), .reg_activation12(reg_activation31_3_1), .reg_activation22(reg_activation31_3_2), .weight_en(weight_en));
SA22 U31_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_4_1), .partial_sum_in12(reg_psum30_4_2), .weight_in11(reg_weight30_4_1), .weight_in12(reg_weight30_4_2), .activation_in11(reg_activation31_3_1), .activation_in21(reg_activation31_3_2), .reg_partial_sum21(reg_psum31_4_1), .reg_partial_sum22(reg_psum31_4_2), .reg_weight21(reg_weight31_4_1), .reg_weight22(reg_weight31_4_2), .reg_activation12(reg_activation31_4_1), .reg_activation22(reg_activation31_4_2), .weight_en(weight_en));
SA22 U31_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_5_1), .partial_sum_in12(reg_psum30_5_2), .weight_in11(reg_weight30_5_1), .weight_in12(reg_weight30_5_2), .activation_in11(reg_activation31_4_1), .activation_in21(reg_activation31_4_2), .reg_partial_sum21(reg_psum31_5_1), .reg_partial_sum22(reg_psum31_5_2), .reg_weight21(reg_weight31_5_1), .reg_weight22(reg_weight31_5_2), .reg_activation12(reg_activation31_5_1), .reg_activation22(reg_activation31_5_2), .weight_en(weight_en));
SA22 U31_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_6_1), .partial_sum_in12(reg_psum30_6_2), .weight_in11(reg_weight30_6_1), .weight_in12(reg_weight30_6_2), .activation_in11(reg_activation31_5_1), .activation_in21(reg_activation31_5_2), .reg_partial_sum21(reg_psum31_6_1), .reg_partial_sum22(reg_psum31_6_2), .reg_weight21(reg_weight31_6_1), .reg_weight22(reg_weight31_6_2), .reg_activation12(reg_activation31_6_1), .reg_activation22(reg_activation31_6_2), .weight_en(weight_en));
SA22 U31_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_7_1), .partial_sum_in12(reg_psum30_7_2), .weight_in11(reg_weight30_7_1), .weight_in12(reg_weight30_7_2), .activation_in11(reg_activation31_6_1), .activation_in21(reg_activation31_6_2), .reg_partial_sum21(reg_psum31_7_1), .reg_partial_sum22(reg_psum31_7_2), .reg_weight21(reg_weight31_7_1), .reg_weight22(reg_weight31_7_2), .reg_activation12(reg_activation31_7_1), .reg_activation22(reg_activation31_7_2), .weight_en(weight_en));
SA22 U31_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_8_1), .partial_sum_in12(reg_psum30_8_2), .weight_in11(reg_weight30_8_1), .weight_in12(reg_weight30_8_2), .activation_in11(reg_activation31_7_1), .activation_in21(reg_activation31_7_2), .reg_partial_sum21(reg_psum31_8_1), .reg_partial_sum22(reg_psum31_8_2), .reg_weight21(reg_weight31_8_1), .reg_weight22(reg_weight31_8_2), .reg_activation12(reg_activation31_8_1), .reg_activation22(reg_activation31_8_2), .weight_en(weight_en));
SA22 U31_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_9_1), .partial_sum_in12(reg_psum30_9_2), .weight_in11(reg_weight30_9_1), .weight_in12(reg_weight30_9_2), .activation_in11(reg_activation31_8_1), .activation_in21(reg_activation31_8_2), .reg_partial_sum21(reg_psum31_9_1), .reg_partial_sum22(reg_psum31_9_2), .reg_weight21(reg_weight31_9_1), .reg_weight22(reg_weight31_9_2), .reg_activation12(reg_activation31_9_1), .reg_activation22(reg_activation31_9_2), .weight_en(weight_en));
SA22 U31_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_10_1), .partial_sum_in12(reg_psum30_10_2), .weight_in11(reg_weight30_10_1), .weight_in12(reg_weight30_10_2), .activation_in11(reg_activation31_9_1), .activation_in21(reg_activation31_9_2), .reg_partial_sum21(reg_psum31_10_1), .reg_partial_sum22(reg_psum31_10_2), .reg_weight21(reg_weight31_10_1), .reg_weight22(reg_weight31_10_2), .reg_activation12(reg_activation31_10_1), .reg_activation22(reg_activation31_10_2), .weight_en(weight_en));
SA22 U31_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_11_1), .partial_sum_in12(reg_psum30_11_2), .weight_in11(reg_weight30_11_1), .weight_in12(reg_weight30_11_2), .activation_in11(reg_activation31_10_1), .activation_in21(reg_activation31_10_2), .reg_partial_sum21(reg_psum31_11_1), .reg_partial_sum22(reg_psum31_11_2), .reg_weight21(reg_weight31_11_1), .reg_weight22(reg_weight31_11_2), .reg_activation12(reg_activation31_11_1), .reg_activation22(reg_activation31_11_2), .weight_en(weight_en));
SA22 U31_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_12_1), .partial_sum_in12(reg_psum30_12_2), .weight_in11(reg_weight30_12_1), .weight_in12(reg_weight30_12_2), .activation_in11(reg_activation31_11_1), .activation_in21(reg_activation31_11_2), .reg_partial_sum21(reg_psum31_12_1), .reg_partial_sum22(reg_psum31_12_2), .reg_weight21(reg_weight31_12_1), .reg_weight22(reg_weight31_12_2), .reg_activation12(reg_activation31_12_1), .reg_activation22(reg_activation31_12_2), .weight_en(weight_en));
SA22 U31_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_13_1), .partial_sum_in12(reg_psum30_13_2), .weight_in11(reg_weight30_13_1), .weight_in12(reg_weight30_13_2), .activation_in11(reg_activation31_12_1), .activation_in21(reg_activation31_12_2), .reg_partial_sum21(reg_psum31_13_1), .reg_partial_sum22(reg_psum31_13_2), .reg_weight21(reg_weight31_13_1), .reg_weight22(reg_weight31_13_2), .reg_activation12(reg_activation31_13_1), .reg_activation22(reg_activation31_13_2), .weight_en(weight_en));
SA22 U31_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_14_1), .partial_sum_in12(reg_psum30_14_2), .weight_in11(reg_weight30_14_1), .weight_in12(reg_weight30_14_2), .activation_in11(reg_activation31_13_1), .activation_in21(reg_activation31_13_2), .reg_partial_sum21(reg_psum31_14_1), .reg_partial_sum22(reg_psum31_14_2), .reg_weight21(reg_weight31_14_1), .reg_weight22(reg_weight31_14_2), .reg_activation12(reg_activation31_14_1), .reg_activation22(reg_activation31_14_2), .weight_en(weight_en));
SA22 U31_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_15_1), .partial_sum_in12(reg_psum30_15_2), .weight_in11(reg_weight30_15_1), .weight_in12(reg_weight30_15_2), .activation_in11(reg_activation31_14_1), .activation_in21(reg_activation31_14_2), .reg_partial_sum21(reg_psum31_15_1), .reg_partial_sum22(reg_psum31_15_2), .reg_weight21(reg_weight31_15_1), .reg_weight22(reg_weight31_15_2), .reg_activation12(reg_activation31_15_1), .reg_activation22(reg_activation31_15_2), .weight_en(weight_en));
SA22 U31_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_16_1), .partial_sum_in12(reg_psum30_16_2), .weight_in11(reg_weight30_16_1), .weight_in12(reg_weight30_16_2), .activation_in11(reg_activation31_15_1), .activation_in21(reg_activation31_15_2), .reg_partial_sum21(reg_psum31_16_1), .reg_partial_sum22(reg_psum31_16_2), .reg_weight21(reg_weight31_16_1), .reg_weight22(reg_weight31_16_2), .reg_activation12(reg_activation31_16_1), .reg_activation22(reg_activation31_16_2), .weight_en(weight_en));
SA22 U31_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_17_1), .partial_sum_in12(reg_psum30_17_2), .weight_in11(reg_weight30_17_1), .weight_in12(reg_weight30_17_2), .activation_in11(reg_activation31_16_1), .activation_in21(reg_activation31_16_2), .reg_partial_sum21(reg_psum31_17_1), .reg_partial_sum22(reg_psum31_17_2), .reg_weight21(reg_weight31_17_1), .reg_weight22(reg_weight31_17_2), .reg_activation12(reg_activation31_17_1), .reg_activation22(reg_activation31_17_2), .weight_en(weight_en));
SA22 U31_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_18_1), .partial_sum_in12(reg_psum30_18_2), .weight_in11(reg_weight30_18_1), .weight_in12(reg_weight30_18_2), .activation_in11(reg_activation31_17_1), .activation_in21(reg_activation31_17_2), .reg_partial_sum21(reg_psum31_18_1), .reg_partial_sum22(reg_psum31_18_2), .reg_weight21(reg_weight31_18_1), .reg_weight22(reg_weight31_18_2), .reg_activation12(reg_activation31_18_1), .reg_activation22(reg_activation31_18_2), .weight_en(weight_en));
SA22 U31_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_19_1), .partial_sum_in12(reg_psum30_19_2), .weight_in11(reg_weight30_19_1), .weight_in12(reg_weight30_19_2), .activation_in11(reg_activation31_18_1), .activation_in21(reg_activation31_18_2), .reg_partial_sum21(reg_psum31_19_1), .reg_partial_sum22(reg_psum31_19_2), .reg_weight21(reg_weight31_19_1), .reg_weight22(reg_weight31_19_2), .reg_activation12(reg_activation31_19_1), .reg_activation22(reg_activation31_19_2), .weight_en(weight_en));
SA22 U31_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_20_1), .partial_sum_in12(reg_psum30_20_2), .weight_in11(reg_weight30_20_1), .weight_in12(reg_weight30_20_2), .activation_in11(reg_activation31_19_1), .activation_in21(reg_activation31_19_2), .reg_partial_sum21(reg_psum31_20_1), .reg_partial_sum22(reg_psum31_20_2), .reg_weight21(reg_weight31_20_1), .reg_weight22(reg_weight31_20_2), .reg_activation12(reg_activation31_20_1), .reg_activation22(reg_activation31_20_2), .weight_en(weight_en));
SA22 U31_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_21_1), .partial_sum_in12(reg_psum30_21_2), .weight_in11(reg_weight30_21_1), .weight_in12(reg_weight30_21_2), .activation_in11(reg_activation31_20_1), .activation_in21(reg_activation31_20_2), .reg_partial_sum21(reg_psum31_21_1), .reg_partial_sum22(reg_psum31_21_2), .reg_weight21(reg_weight31_21_1), .reg_weight22(reg_weight31_21_2), .reg_activation12(reg_activation31_21_1), .reg_activation22(reg_activation31_21_2), .weight_en(weight_en));
SA22 U31_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_22_1), .partial_sum_in12(reg_psum30_22_2), .weight_in11(reg_weight30_22_1), .weight_in12(reg_weight30_22_2), .activation_in11(reg_activation31_21_1), .activation_in21(reg_activation31_21_2), .reg_partial_sum21(reg_psum31_22_1), .reg_partial_sum22(reg_psum31_22_2), .reg_weight21(reg_weight31_22_1), .reg_weight22(reg_weight31_22_2), .reg_activation12(reg_activation31_22_1), .reg_activation22(reg_activation31_22_2), .weight_en(weight_en));
SA22 U31_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_23_1), .partial_sum_in12(reg_psum30_23_2), .weight_in11(reg_weight30_23_1), .weight_in12(reg_weight30_23_2), .activation_in11(reg_activation31_22_1), .activation_in21(reg_activation31_22_2), .reg_partial_sum21(reg_psum31_23_1), .reg_partial_sum22(reg_psum31_23_2), .reg_weight21(reg_weight31_23_1), .reg_weight22(reg_weight31_23_2), .reg_activation12(reg_activation31_23_1), .reg_activation22(reg_activation31_23_2), .weight_en(weight_en));
SA22 U31_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_24_1), .partial_sum_in12(reg_psum30_24_2), .weight_in11(reg_weight30_24_1), .weight_in12(reg_weight30_24_2), .activation_in11(reg_activation31_23_1), .activation_in21(reg_activation31_23_2), .reg_partial_sum21(reg_psum31_24_1), .reg_partial_sum22(reg_psum31_24_2), .reg_weight21(reg_weight31_24_1), .reg_weight22(reg_weight31_24_2), .reg_activation12(reg_activation31_24_1), .reg_activation22(reg_activation31_24_2), .weight_en(weight_en));
SA22 U31_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_25_1), .partial_sum_in12(reg_psum30_25_2), .weight_in11(reg_weight30_25_1), .weight_in12(reg_weight30_25_2), .activation_in11(reg_activation31_24_1), .activation_in21(reg_activation31_24_2), .reg_partial_sum21(reg_psum31_25_1), .reg_partial_sum22(reg_psum31_25_2), .reg_weight21(reg_weight31_25_1), .reg_weight22(reg_weight31_25_2), .reg_activation12(reg_activation31_25_1), .reg_activation22(reg_activation31_25_2), .weight_en(weight_en));
SA22 U31_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_26_1), .partial_sum_in12(reg_psum30_26_2), .weight_in11(reg_weight30_26_1), .weight_in12(reg_weight30_26_2), .activation_in11(reg_activation31_25_1), .activation_in21(reg_activation31_25_2), .reg_partial_sum21(reg_psum31_26_1), .reg_partial_sum22(reg_psum31_26_2), .reg_weight21(reg_weight31_26_1), .reg_weight22(reg_weight31_26_2), .reg_activation12(reg_activation31_26_1), .reg_activation22(reg_activation31_26_2), .weight_en(weight_en));
SA22 U31_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_27_1), .partial_sum_in12(reg_psum30_27_2), .weight_in11(reg_weight30_27_1), .weight_in12(reg_weight30_27_2), .activation_in11(reg_activation31_26_1), .activation_in21(reg_activation31_26_2), .reg_partial_sum21(reg_psum31_27_1), .reg_partial_sum22(reg_psum31_27_2), .reg_weight21(reg_weight31_27_1), .reg_weight22(reg_weight31_27_2), .reg_activation12(reg_activation31_27_1), .reg_activation22(reg_activation31_27_2), .weight_en(weight_en));
SA22 U31_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_28_1), .partial_sum_in12(reg_psum30_28_2), .weight_in11(reg_weight30_28_1), .weight_in12(reg_weight30_28_2), .activation_in11(reg_activation31_27_1), .activation_in21(reg_activation31_27_2), .reg_partial_sum21(reg_psum31_28_1), .reg_partial_sum22(reg_psum31_28_2), .reg_weight21(reg_weight31_28_1), .reg_weight22(reg_weight31_28_2), .reg_activation12(reg_activation31_28_1), .reg_activation22(reg_activation31_28_2), .weight_en(weight_en));
SA22 U31_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_29_1), .partial_sum_in12(reg_psum30_29_2), .weight_in11(reg_weight30_29_1), .weight_in12(reg_weight30_29_2), .activation_in11(reg_activation31_28_1), .activation_in21(reg_activation31_28_2), .reg_partial_sum21(reg_psum31_29_1), .reg_partial_sum22(reg_psum31_29_2), .reg_weight21(reg_weight31_29_1), .reg_weight22(reg_weight31_29_2), .reg_activation12(reg_activation31_29_1), .reg_activation22(reg_activation31_29_2), .weight_en(weight_en));
SA22 U31_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_30_1), .partial_sum_in12(reg_psum30_30_2), .weight_in11(reg_weight30_30_1), .weight_in12(reg_weight30_30_2), .activation_in11(reg_activation31_29_1), .activation_in21(reg_activation31_29_2), .reg_partial_sum21(reg_psum31_30_1), .reg_partial_sum22(reg_psum31_30_2), .reg_weight21(reg_weight31_30_1), .reg_weight22(reg_weight31_30_2), .reg_activation12(reg_activation31_30_1), .reg_activation22(reg_activation31_30_2), .weight_en(weight_en));
SA22 U31_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_31_1), .partial_sum_in12(reg_psum30_31_2), .weight_in11(reg_weight30_31_1), .weight_in12(reg_weight30_31_2), .activation_in11(reg_activation31_30_1), .activation_in21(reg_activation31_30_2), .reg_partial_sum21(reg_psum31_31_1), .reg_partial_sum22(reg_psum31_31_2), .reg_weight21(reg_weight31_31_1), .reg_weight22(reg_weight31_31_2), .reg_activation12(reg_activation31_31_1), .reg_activation22(reg_activation31_31_2), .weight_en(weight_en));
SA22 U31_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum30_32_1), .partial_sum_in12(reg_psum30_32_2), .weight_in11(reg_weight30_32_1), .weight_in12(reg_weight30_32_2), .activation_in11(reg_activation31_31_1), .activation_in21(reg_activation31_31_2), .reg_partial_sum21(reg_psum31_32_1), .reg_partial_sum22(reg_psum31_32_2), .reg_weight21(reg_weight31_32_1), .reg_weight22(reg_weight31_32_2), .weight_en(weight_en));
SA22 U32_1(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_1_1), .partial_sum_in12(reg_psum31_1_2), .weight_in11(reg_weight31_1_1), .weight_in12(reg_weight31_1_2), .activation_in11(in_activation32_1_1), .activation_in21(in_activation32_1_2), .reg_partial_sum21(reg_psum32_1_1), .reg_partial_sum22(reg_psum32_1_2), .reg_activation12(reg_activation32_1_1), .reg_activation22(reg_activation32_1_2), .weight_en(weight_en));
SA22 U32_2(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_2_1), .partial_sum_in12(reg_psum31_2_2), .weight_in11(reg_weight31_2_1), .weight_in12(reg_weight31_2_2), .activation_in11(reg_activation32_1_1), .activation_in21(reg_activation32_1_2), .reg_partial_sum21(reg_psum32_2_1), .reg_partial_sum22(reg_psum32_2_2), .reg_activation12(reg_activation32_2_1), .reg_activation22(reg_activation32_2_2), .weight_en(weight_en));
SA22 U32_3(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_3_1), .partial_sum_in12(reg_psum31_3_2), .weight_in11(reg_weight31_3_1), .weight_in12(reg_weight31_3_2), .activation_in11(reg_activation32_2_1), .activation_in21(reg_activation32_2_2), .reg_partial_sum21(reg_psum32_3_1), .reg_partial_sum22(reg_psum32_3_2), .reg_activation12(reg_activation32_3_1), .reg_activation22(reg_activation32_3_2), .weight_en(weight_en));
SA22 U32_4(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_4_1), .partial_sum_in12(reg_psum31_4_2), .weight_in11(reg_weight31_4_1), .weight_in12(reg_weight31_4_2), .activation_in11(reg_activation32_3_1), .activation_in21(reg_activation32_3_2), .reg_partial_sum21(reg_psum32_4_1), .reg_partial_sum22(reg_psum32_4_2), .reg_activation12(reg_activation32_4_1), .reg_activation22(reg_activation32_4_2), .weight_en(weight_en));
SA22 U32_5(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_5_1), .partial_sum_in12(reg_psum31_5_2), .weight_in11(reg_weight31_5_1), .weight_in12(reg_weight31_5_2), .activation_in11(reg_activation32_4_1), .activation_in21(reg_activation32_4_2), .reg_partial_sum21(reg_psum32_5_1), .reg_partial_sum22(reg_psum32_5_2), .reg_activation12(reg_activation32_5_1), .reg_activation22(reg_activation32_5_2), .weight_en(weight_en));
SA22 U32_6(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_6_1), .partial_sum_in12(reg_psum31_6_2), .weight_in11(reg_weight31_6_1), .weight_in12(reg_weight31_6_2), .activation_in11(reg_activation32_5_1), .activation_in21(reg_activation32_5_2), .reg_partial_sum21(reg_psum32_6_1), .reg_partial_sum22(reg_psum32_6_2), .reg_activation12(reg_activation32_6_1), .reg_activation22(reg_activation32_6_2), .weight_en(weight_en));
SA22 U32_7(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_7_1), .partial_sum_in12(reg_psum31_7_2), .weight_in11(reg_weight31_7_1), .weight_in12(reg_weight31_7_2), .activation_in11(reg_activation32_6_1), .activation_in21(reg_activation32_6_2), .reg_partial_sum21(reg_psum32_7_1), .reg_partial_sum22(reg_psum32_7_2), .reg_activation12(reg_activation32_7_1), .reg_activation22(reg_activation32_7_2), .weight_en(weight_en));
SA22 U32_8(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_8_1), .partial_sum_in12(reg_psum31_8_2), .weight_in11(reg_weight31_8_1), .weight_in12(reg_weight31_8_2), .activation_in11(reg_activation32_7_1), .activation_in21(reg_activation32_7_2), .reg_partial_sum21(reg_psum32_8_1), .reg_partial_sum22(reg_psum32_8_2), .reg_activation12(reg_activation32_8_1), .reg_activation22(reg_activation32_8_2), .weight_en(weight_en));
SA22 U32_9(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_9_1), .partial_sum_in12(reg_psum31_9_2), .weight_in11(reg_weight31_9_1), .weight_in12(reg_weight31_9_2), .activation_in11(reg_activation32_8_1), .activation_in21(reg_activation32_8_2), .reg_partial_sum21(reg_psum32_9_1), .reg_partial_sum22(reg_psum32_9_2), .reg_activation12(reg_activation32_9_1), .reg_activation22(reg_activation32_9_2), .weight_en(weight_en));
SA22 U32_10(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_10_1), .partial_sum_in12(reg_psum31_10_2), .weight_in11(reg_weight31_10_1), .weight_in12(reg_weight31_10_2), .activation_in11(reg_activation32_9_1), .activation_in21(reg_activation32_9_2), .reg_partial_sum21(reg_psum32_10_1), .reg_partial_sum22(reg_psum32_10_2), .reg_activation12(reg_activation32_10_1), .reg_activation22(reg_activation32_10_2), .weight_en(weight_en));
SA22 U32_11(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_11_1), .partial_sum_in12(reg_psum31_11_2), .weight_in11(reg_weight31_11_1), .weight_in12(reg_weight31_11_2), .activation_in11(reg_activation32_10_1), .activation_in21(reg_activation32_10_2), .reg_partial_sum21(reg_psum32_11_1), .reg_partial_sum22(reg_psum32_11_2), .reg_activation12(reg_activation32_11_1), .reg_activation22(reg_activation32_11_2), .weight_en(weight_en));
SA22 U32_12(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_12_1), .partial_sum_in12(reg_psum31_12_2), .weight_in11(reg_weight31_12_1), .weight_in12(reg_weight31_12_2), .activation_in11(reg_activation32_11_1), .activation_in21(reg_activation32_11_2), .reg_partial_sum21(reg_psum32_12_1), .reg_partial_sum22(reg_psum32_12_2), .reg_activation12(reg_activation32_12_1), .reg_activation22(reg_activation32_12_2), .weight_en(weight_en));
SA22 U32_13(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_13_1), .partial_sum_in12(reg_psum31_13_2), .weight_in11(reg_weight31_13_1), .weight_in12(reg_weight31_13_2), .activation_in11(reg_activation32_12_1), .activation_in21(reg_activation32_12_2), .reg_partial_sum21(reg_psum32_13_1), .reg_partial_sum22(reg_psum32_13_2), .reg_activation12(reg_activation32_13_1), .reg_activation22(reg_activation32_13_2), .weight_en(weight_en));
SA22 U32_14(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_14_1), .partial_sum_in12(reg_psum31_14_2), .weight_in11(reg_weight31_14_1), .weight_in12(reg_weight31_14_2), .activation_in11(reg_activation32_13_1), .activation_in21(reg_activation32_13_2), .reg_partial_sum21(reg_psum32_14_1), .reg_partial_sum22(reg_psum32_14_2), .reg_activation12(reg_activation32_14_1), .reg_activation22(reg_activation32_14_2), .weight_en(weight_en));
SA22 U32_15(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_15_1), .partial_sum_in12(reg_psum31_15_2), .weight_in11(reg_weight31_15_1), .weight_in12(reg_weight31_15_2), .activation_in11(reg_activation32_14_1), .activation_in21(reg_activation32_14_2), .reg_partial_sum21(reg_psum32_15_1), .reg_partial_sum22(reg_psum32_15_2), .reg_activation12(reg_activation32_15_1), .reg_activation22(reg_activation32_15_2), .weight_en(weight_en));
SA22 U32_16(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_16_1), .partial_sum_in12(reg_psum31_16_2), .weight_in11(reg_weight31_16_1), .weight_in12(reg_weight31_16_2), .activation_in11(reg_activation32_15_1), .activation_in21(reg_activation32_15_2), .reg_partial_sum21(reg_psum32_16_1), .reg_partial_sum22(reg_psum32_16_2), .reg_activation12(reg_activation32_16_1), .reg_activation22(reg_activation32_16_2), .weight_en(weight_en));
SA22 U32_17(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_17_1), .partial_sum_in12(reg_psum31_17_2), .weight_in11(reg_weight31_17_1), .weight_in12(reg_weight31_17_2), .activation_in11(reg_activation32_16_1), .activation_in21(reg_activation32_16_2), .reg_partial_sum21(reg_psum32_17_1), .reg_partial_sum22(reg_psum32_17_2), .reg_activation12(reg_activation32_17_1), .reg_activation22(reg_activation32_17_2), .weight_en(weight_en));
SA22 U32_18(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_18_1), .partial_sum_in12(reg_psum31_18_2), .weight_in11(reg_weight31_18_1), .weight_in12(reg_weight31_18_2), .activation_in11(reg_activation32_17_1), .activation_in21(reg_activation32_17_2), .reg_partial_sum21(reg_psum32_18_1), .reg_partial_sum22(reg_psum32_18_2), .reg_activation12(reg_activation32_18_1), .reg_activation22(reg_activation32_18_2), .weight_en(weight_en));
SA22 U32_19(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_19_1), .partial_sum_in12(reg_psum31_19_2), .weight_in11(reg_weight31_19_1), .weight_in12(reg_weight31_19_2), .activation_in11(reg_activation32_18_1), .activation_in21(reg_activation32_18_2), .reg_partial_sum21(reg_psum32_19_1), .reg_partial_sum22(reg_psum32_19_2), .reg_activation12(reg_activation32_19_1), .reg_activation22(reg_activation32_19_2), .weight_en(weight_en));
SA22 U32_20(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_20_1), .partial_sum_in12(reg_psum31_20_2), .weight_in11(reg_weight31_20_1), .weight_in12(reg_weight31_20_2), .activation_in11(reg_activation32_19_1), .activation_in21(reg_activation32_19_2), .reg_partial_sum21(reg_psum32_20_1), .reg_partial_sum22(reg_psum32_20_2), .reg_activation12(reg_activation32_20_1), .reg_activation22(reg_activation32_20_2), .weight_en(weight_en));
SA22 U32_21(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_21_1), .partial_sum_in12(reg_psum31_21_2), .weight_in11(reg_weight31_21_1), .weight_in12(reg_weight31_21_2), .activation_in11(reg_activation32_20_1), .activation_in21(reg_activation32_20_2), .reg_partial_sum21(reg_psum32_21_1), .reg_partial_sum22(reg_psum32_21_2), .reg_activation12(reg_activation32_21_1), .reg_activation22(reg_activation32_21_2), .weight_en(weight_en));
SA22 U32_22(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_22_1), .partial_sum_in12(reg_psum31_22_2), .weight_in11(reg_weight31_22_1), .weight_in12(reg_weight31_22_2), .activation_in11(reg_activation32_21_1), .activation_in21(reg_activation32_21_2), .reg_partial_sum21(reg_psum32_22_1), .reg_partial_sum22(reg_psum32_22_2), .reg_activation12(reg_activation32_22_1), .reg_activation22(reg_activation32_22_2), .weight_en(weight_en));
SA22 U32_23(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_23_1), .partial_sum_in12(reg_psum31_23_2), .weight_in11(reg_weight31_23_1), .weight_in12(reg_weight31_23_2), .activation_in11(reg_activation32_22_1), .activation_in21(reg_activation32_22_2), .reg_partial_sum21(reg_psum32_23_1), .reg_partial_sum22(reg_psum32_23_2), .reg_activation12(reg_activation32_23_1), .reg_activation22(reg_activation32_23_2), .weight_en(weight_en));
SA22 U32_24(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_24_1), .partial_sum_in12(reg_psum31_24_2), .weight_in11(reg_weight31_24_1), .weight_in12(reg_weight31_24_2), .activation_in11(reg_activation32_23_1), .activation_in21(reg_activation32_23_2), .reg_partial_sum21(reg_psum32_24_1), .reg_partial_sum22(reg_psum32_24_2), .reg_activation12(reg_activation32_24_1), .reg_activation22(reg_activation32_24_2), .weight_en(weight_en));
SA22 U32_25(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_25_1), .partial_sum_in12(reg_psum31_25_2), .weight_in11(reg_weight31_25_1), .weight_in12(reg_weight31_25_2), .activation_in11(reg_activation32_24_1), .activation_in21(reg_activation32_24_2), .reg_partial_sum21(reg_psum32_25_1), .reg_partial_sum22(reg_psum32_25_2), .reg_activation12(reg_activation32_25_1), .reg_activation22(reg_activation32_25_2), .weight_en(weight_en));
SA22 U32_26(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_26_1), .partial_sum_in12(reg_psum31_26_2), .weight_in11(reg_weight31_26_1), .weight_in12(reg_weight31_26_2), .activation_in11(reg_activation32_25_1), .activation_in21(reg_activation32_25_2), .reg_partial_sum21(reg_psum32_26_1), .reg_partial_sum22(reg_psum32_26_2), .reg_activation12(reg_activation32_26_1), .reg_activation22(reg_activation32_26_2), .weight_en(weight_en));
SA22 U32_27(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_27_1), .partial_sum_in12(reg_psum31_27_2), .weight_in11(reg_weight31_27_1), .weight_in12(reg_weight31_27_2), .activation_in11(reg_activation32_26_1), .activation_in21(reg_activation32_26_2), .reg_partial_sum21(reg_psum32_27_1), .reg_partial_sum22(reg_psum32_27_2), .reg_activation12(reg_activation32_27_1), .reg_activation22(reg_activation32_27_2), .weight_en(weight_en));
SA22 U32_28(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_28_1), .partial_sum_in12(reg_psum31_28_2), .weight_in11(reg_weight31_28_1), .weight_in12(reg_weight31_28_2), .activation_in11(reg_activation32_27_1), .activation_in21(reg_activation32_27_2), .reg_partial_sum21(reg_psum32_28_1), .reg_partial_sum22(reg_psum32_28_2), .reg_activation12(reg_activation32_28_1), .reg_activation22(reg_activation32_28_2), .weight_en(weight_en));
SA22 U32_29(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_29_1), .partial_sum_in12(reg_psum31_29_2), .weight_in11(reg_weight31_29_1), .weight_in12(reg_weight31_29_2), .activation_in11(reg_activation32_28_1), .activation_in21(reg_activation32_28_2), .reg_partial_sum21(reg_psum32_29_1), .reg_partial_sum22(reg_psum32_29_2), .reg_activation12(reg_activation32_29_1), .reg_activation22(reg_activation32_29_2), .weight_en(weight_en));
SA22 U32_30(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_30_1), .partial_sum_in12(reg_psum31_30_2), .weight_in11(reg_weight31_30_1), .weight_in12(reg_weight31_30_2), .activation_in11(reg_activation32_29_1), .activation_in21(reg_activation32_29_2), .reg_partial_sum21(reg_psum32_30_1), .reg_partial_sum22(reg_psum32_30_2), .reg_activation12(reg_activation32_30_1), .reg_activation22(reg_activation32_30_2), .weight_en(weight_en));
SA22 U32_31(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_31_1), .partial_sum_in12(reg_psum31_31_2), .weight_in11(reg_weight31_31_1), .weight_in12(reg_weight31_31_2), .activation_in11(reg_activation32_30_1), .activation_in21(reg_activation32_30_2), .reg_partial_sum21(reg_psum32_31_1), .reg_partial_sum22(reg_psum32_31_2), .reg_activation12(reg_activation32_31_1), .reg_activation22(reg_activation32_31_2), .weight_en(weight_en));
SA22 U32_32(.clk(clk), .rst(rst), .partial_sum_in11(reg_psum31_32_1), .partial_sum_in12(reg_psum31_32_2), .weight_in11(reg_weight31_32_1), .weight_in12(reg_weight31_32_2), .activation_in11(reg_activation32_31_1), .activation_in21(reg_activation32_31_2), .reg_partial_sum21(reg_psum32_32_1), .reg_partial_sum22(reg_psum32_32_2), .weight_en(weight_en));
endmodule